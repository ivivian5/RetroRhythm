library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity arrow_rom is 
 	port(
		outglobal_o : in std_logic;
		addr_x : in std_logic_vector(4 downto 0);
		addr_y : in std_logic_vector(4 downto 0);
		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
	);
end;

architecture sim of arrow_rom is
signal addr : std_logic_vector(9 downto 0);

begin
	addr (9 downto 5) <= addr_y;
	addr (4 downto 0) <= addr_x;
	process(outglobal_o) begin
		if rising_edge(outglobal_o) then
			case addr is
				when "0000000111" => data <= "110011";
				when "0000100110" => data <= "110011";
				when "0000100111" => data <= "110011";
				when "0000101000" => data <= "110011";
				when "0001000101" => data <= "110011";
				when "0001000110" => data <= "110011";
				when "0001000111" => data <= "111111";
				when "0001001000" => data <= "110011";
				when "0001100100" => data <= "110011";
				when "0001100101" => data <= "110011";
				when "0001100110" => data <= "111111";
				when "0001100111" => data <= "110011";
				when "0001101000" => data <= "110011";
				when "0010000011" => data <= "110011";
				when "0010000100" => data <= "110011";
				when "0010000101" => data <= "111111";
				when "0010000110" => data <= "110011";
				when "0010000111" => data <= "110011";
				when "0010001000" => data <= "110011";
				when "0010100010" => data <= "110011";
				when "0010100011" => data <= "110011";
				when "0010100100" => data <= "111111";
				when "0010100101" => data <= "110011";
				when "0010100110" => data <= "110011";
				when "0010100111" => data <= "110011";
				when "0010101000" => data <= "110011";
				when "0010101001" => data <= "110011";
				when "0010101010" => data <= "110011";
				when "0010101011" => data <= "110011";
				when "0010101100" => data <= "110011";
				when "0010101101" => data <= "110011";
				when "0011000001" => data <= "110011";
				when "0011000010" => data <= "110011";
				when "0011000011" => data <= "111111";
				when "0011000100" => data <= "110011";
				when "0011000101" => data <= "110011";
				when "0011000110" => data <= "110011";
				when "0011000111" => data <= "110011";
				when "0011001000" => data <= "110011";
				when "0011001001" => data <= "110011";
				when "0011001010" => data <= "110011";
				when "0011001011" => data <= "110011";
				when "0011001100" => data <= "110011";
				when "0011001101" => data <= "110011";
				when "0011001110" => data <= "110011";
				when "0011100000" => data <= "110011";
				when "0011100001" => data <= "110011";
				when "0011100010" => data <= "111111";
				when "0011100011" => data <= "110011";
				when "0011100100" => data <= "110011";
				when "0011100101" => data <= "110011";
				when "0011100110" => data <= "110011";
				when "0011100111" => data <= "110011";
				when "0011101000" => data <= "110011";
				when "0011101001" => data <= "110011";
				when "0011101010" => data <= "110011";
				when "0011101011" => data <= "110011";
				when "0011101100" => data <= "110011";
				when "0011101101" => data <= "110011";
				when "0011101110" => data <= "110011";
				when "0100000001" => data <= "110011";
				when "0100000010" => data <= "110011";
				when "0100000011" => data <= "110011";
				when "0100000100" => data <= "110011";
				when "0100000101" => data <= "110011";
				when "0100000110" => data <= "110011";
				when "0100000111" => data <= "110011";
				when "0100001000" => data <= "110011";
				when "0100001001" => data <= "110011";
				when "0100001010" => data <= "110011";
				when "0100001011" => data <= "110011";
				when "0100001100" => data <= "110011";
				when "0100001101" => data <= "110011";
				when "0100001110" => data <= "110011";
				when "0100100010" => data <= "110011";
				when "0100100011" => data <= "110011";
				when "0100100100" => data <= "110011";
				when "0100100101" => data <= "110011";
				when "0100100110" => data <= "110011";
				when "0100100111" => data <= "110011";
				when "0100101000" => data <= "110011";
				when "0100101001" => data <= "110011";
				when "0100101010" => data <= "110011";
				when "0100101011" => data <= "110011";
				when "0100101100" => data <= "110011";
				when "0100101101" => data <= "110011";
				when "0101000011" => data <= "110011";
				when "0101000100" => data <= "110011";
				when "0101000101" => data <= "110011";
				when "0101000110" => data <= "110011";
				when "0101000111" => data <= "110011";
				when "0101001000" => data <= "110011";
				when "0101100100" => data <= "110011";
				when "0101100101" => data <= "110011";
				when "0101100110" => data <= "110011";
				when "0101100111" => data <= "110011";
				when "0101101000" => data <= "110011";
				when "0110000101" => data <= "110011";
				when "0110000110" => data <= "110011";
				when "0110000111" => data <= "110011";
				when "0110001000" => data <= "110011";
				when "0110100110" => data <= "110011";
				when "0110100111" => data <= "110011";
				when "0110101000" => data <= "110011";
				when "0111000111" => data <= "110011";
				when others => data <= "000001";
			end case;
		end if; 
	end process; 
end;