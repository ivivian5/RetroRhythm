library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity rom is
                	port(
                		clk : in std_logic;
                		addr : in std_logic_vector(3 downto 0); -- 16 words total
                		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
                	);
                end;

                architecture sim of rom is
                begin
                	process(clk) begin
                		if rising_edge(clk) then
                			case addr is
				when "000000000000" => data <= "000000";
				when "000000000001" => data <= "000000";
				when "000000000010" => data <= "000000";
				when "000000000011" => data <= "000000";
				when "000000000100" => data <= "000000";
				when "000000000101" => data <= "000000";
				when "000000000110" => data <= "000000";
				when "000000000111" => data <= "000000";
				when "000000001000" => data <= "000000";
				when "000000001001" => data <= "000000";
				when "000000001010" => data <= "000000";
				when "000000001011" => data <= "000000";
				when "000000001100" => data <= "000000";
				when "000000001101" => data <= "000000";
				when "000000001110" => data <= "000000";
				when "000000001111" => data <= "000000";
				when "000000010000" => data <= "000000";
				when "000000010001" => data <= "000000";
				when "000000010010" => data <= "000000";
				when "000000010011" => data <= "000000";
				when "000000010100" => data <= "000000";
				when "000000010101" => data <= "000000";
				when "000000010110" => data <= "000000";
				when "000000010111" => data <= "000000";
				when "000000011000" => data <= "000000";
				when "000000011001" => data <= "000000";
				when "000000011010" => data <= "000000";
				when "000000011011" => data <= "000000";
				when "000000011100" => data <= "000000";
				when "000000011101" => data <= "000000";
				when "000000011110" => data <= "000000";
				when "000000011111" => data <= "000000";
				when "000000100000" => data <= "000000";
				when "000000100001" => data <= "000000";
				when "000000100010" => data <= "000000";
				when "000000100011" => data <= "000000";
				when "000000100100" => data <= "000000";
				when "000000100101" => data <= "000000";
				when "000000100110" => data <= "000000";
				when "000000100111" => data <= "000000";
				when "000000101000" => data <= "000000";
				when "000000101001" => data <= "000000";
				when "000000101010" => data <= "000000";
				when "000000101011" => data <= "000000";
				when "000000101100" => data <= "000000";
				when "000000101101" => data <= "000000";
				when "000000101110" => data <= "000000";
				when "000000101111" => data <= "000000";
				when "000000110000" => data <= "000000";
				when "000000110001" => data <= "000000";
				when "000000110010" => data <= "000000";
				when "000000110011" => data <= "000000";
				when "000000110100" => data <= "000000";
				when "000000110101" => data <= "000000";
				when "000000110110" => data <= "000000";
				when "000000110111" => data <= "000000";
				when "000000111000" => data <= "000000";
				when "000000111001" => data <= "000000";
				when "000000111010" => data <= "000000";
				when "000000111011" => data <= "000000";
				when "000000111100" => data <= "000000";
				when "000000111101" => data <= "000000";
				when "000000111110" => data <= "000000";
				when "000000111111" => data <= "000000";
				when "000001000000" => data <= "000000";
				when "000001000001" => data <= "000000";
				when "000001000010" => data <= "000000";
				when "000001000011" => data <= "000000";
				when "000001000100" => data <= "000000";
				when "000001000101" => data <= "000000";
				when "000001000110" => data <= "000000";
				when "000001000111" => data <= "000000";
				when "000001001000" => data <= "000000";
				when "000001001001" => data <= "000000";
				when "000001001010" => data <= "000000";
				when "000001001011" => data <= "000000";
				when "000001001100" => data <= "000000";
				when "000001001101" => data <= "000000";
				when "000001001110" => data <= "000000";
				when "000001001111" => data <= "000000";
				when "000001010000" => data <= "000000";
				when "000001010001" => data <= "000000";
				when "000001010010" => data <= "000000";
				when "000001010011" => data <= "000000";
				when "000001010100" => data <= "000000";
				when "000001010101" => data <= "000000";
				when "000001010110" => data <= "000000";
				when "000001010111" => data <= "000000";
				when "000001011000" => data <= "000000";
				when "000001011001" => data <= "000000";
				when "000001011010" => data <= "000000";
				when "000001011011" => data <= "000000";
				when "000001011100" => data <= "000000";
				when "000001011101" => data <= "000000";
				when "000001011110" => data <= "000000";
				when "000001011111" => data <= "000000";
				when "000001100000" => data <= "000000";
				when "000001100001" => data <= "000000";
				when "000001100010" => data <= "000000";
				when "000001100011" => data <= "000000";
				when "000001100100" => data <= "000000";
				when "000001100101" => data <= "000000";
				when "000001100110" => data <= "000000";
				when "000001100111" => data <= "000000";
				when "000001101000" => data <= "000000";
				when "000001101001" => data <= "000000";
				when "000001101010" => data <= "000000";
				when "000001101011" => data <= "000000";
				when "000001101100" => data <= "000000";
				when "000001101101" => data <= "000000";
				when "000001101110" => data <= "000000";
				when "000001101111" => data <= "000000";
				when "000001110000" => data <= "000000";
				when "000001110001" => data <= "000000";
				when "000001110010" => data <= "000000";
				when "000001110011" => data <= "000000";
				when "000001110100" => data <= "000000";
				when "000001110101" => data <= "000000";
				when "000001110110" => data <= "000000";
				when "000001110111" => data <= "000000";
				when "000001111000" => data <= "000000";
				when "000001111001" => data <= "000000";
				when "000001111010" => data <= "000000";
				when "000001111011" => data <= "000000";
				when "000001111100" => data <= "000000";
				when "000001111101" => data <= "000000";
				when "000001111110" => data <= "000000";
				when "000001111111" => data <= "000000";
				when "000010000000" => data <= "000000";
				when "000010000001" => data <= "000000";
				when "000010000010" => data <= "000000";
				when "000010000011" => data <= "000000";
				when "000010000100" => data <= "000000";
				when "000010000101" => data <= "000000";
				when "000010000110" => data <= "000000";
				when "000010000111" => data <= "000000";
				when "000010001000" => data <= "000000";
				when "000010001001" => data <= "000000";
				when "000010001010" => data <= "000000";
				when "000010001011" => data <= "000000";
				when "000010001100" => data <= "000000";
				when "000010001101" => data <= "000000";
				when "000010001110" => data <= "000000";
				when "000010001111" => data <= "000000";
				when "000010010000" => data <= "000000";
				when "000010010001" => data <= "000000";
				when "000010010010" => data <= "000000";
				when "000010010011" => data <= "000000";
				when "000010010100" => data <= "000000";
				when "000010010101" => data <= "000000";
				when "000010010110" => data <= "000000";
				when "000010010111" => data <= "000000";
				when "000010011000" => data <= "000000";
				when "000010011001" => data <= "000000";
				when "000010011010" => data <= "000000";
				when "000010011011" => data <= "000000";
				when "000010011100" => data <= "000000";
				when "000010011101" => data <= "000000";
				when "000010011110" => data <= "000000";
				when "000010011111" => data <= "000000";
				when "000010100000" => data <= "000000";
				when "000010100001" => data <= "000000";
				when "000010100010" => data <= "000000";
				when "000010100011" => data <= "000000";
				when "000010100100" => data <= "000000";
				when "000010100101" => data <= "000000";
				when "000010100110" => data <= "000000";
				when "000010100111" => data <= "000000";
				when "000010101000" => data <= "000000";
				when "000010101001" => data <= "000000";
				when "000010101010" => data <= "000000";
				when "000010101011" => data <= "000000";
				when "000010101100" => data <= "000000";
				when "000010101101" => data <= "000000";
				when "000010101110" => data <= "000000";
				when "000010101111" => data <= "000000";
				when "000010110000" => data <= "000000";
				when "000010110001" => data <= "000000";
				when "000010110010" => data <= "000000";
				when "000010110011" => data <= "000000";
				when "000010110100" => data <= "000000";
				when "000010110101" => data <= "000000";
				when "000010110110" => data <= "000000";
				when "000010110111" => data <= "000000";
				when "000010111000" => data <= "000000";
				when "000010111001" => data <= "000000";
				when "000010111010" => data <= "000000";
				when "000010111011" => data <= "000000";
				when "000010111100" => data <= "000000";
				when "000010111101" => data <= "000000";
				when "000010111110" => data <= "000000";
				when "000010111111" => data <= "000000";
				when "000011000000" => data <= "000000";
				when "000011000001" => data <= "000000";
				when "000011000010" => data <= "000000";
				when "000011000011" => data <= "000000";
				when "000011000100" => data <= "000000";
				when "000011000101" => data <= "000000";
				when "000011000110" => data <= "000000";
				when "000011000111" => data <= "000000";
				when "000011001000" => data <= "000000";
				when "000011001001" => data <= "000000";
				when "000011001010" => data <= "000000";
				when "000011001011" => data <= "000000";
				when "000011001100" => data <= "000000";
				when "000011001101" => data <= "000000";
				when "000011001110" => data <= "000000";
				when "000011001111" => data <= "000000";
				when "000011010000" => data <= "000000";
				when "000011010001" => data <= "000000";
				when "000011010010" => data <= "000000";
				when "000011010011" => data <= "000000";
				when "000011010100" => data <= "000000";
				when "000011010101" => data <= "000000";
				when "000011010110" => data <= "000000";
				when "000011010111" => data <= "000000";
				when "000011011000" => data <= "000000";
				when "000011011001" => data <= "000000";
				when "000011011010" => data <= "000000";
				when "000011011011" => data <= "000000";
				when "000011011100" => data <= "000000";
				when "000011011101" => data <= "000000";
				when "000011011110" => data <= "000000";
				when "000011011111" => data <= "000000";
				when "000011100000" => data <= "000000";
				when "000011100001" => data <= "000000";
				when "000011100010" => data <= "000000";
				when "000011100011" => data <= "000000";
				when "000011100100" => data <= "000000";
				when "000011100101" => data <= "000000";
				when "000011100110" => data <= "000000";
				when "000011100111" => data <= "000000";
				when "000011101000" => data <= "000000";
				when "000011101001" => data <= "000000";
				when "000011101010" => data <= "000000";
				when "000011101011" => data <= "000000";
				when "000011101100" => data <= "000000";
				when "000011101101" => data <= "000000";
				when "000011101110" => data <= "000000";
				when "000011101111" => data <= "000000";
				when "000011110000" => data <= "000000";
				when "000011110001" => data <= "000000";
				when "000011110010" => data <= "000000";
				when "000011110011" => data <= "000000";
				when "000011110100" => data <= "000000";
				when "000011110101" => data <= "000000";
				when "000011110110" => data <= "000000";
				when "000011110111" => data <= "000000";
				when "000011111000" => data <= "000000";
				when "000011111001" => data <= "000000";
				when "000011111010" => data <= "000000";
				when "000011111011" => data <= "000000";
				when "000011111100" => data <= "000000";
				when "000011111101" => data <= "000000";
				when "000011111110" => data <= "000000";
				when "000011111111" => data <= "000000";
				when "000100000000" => data <= "000000";
				when "000100000001" => data <= "000000";
				when "000100000010" => data <= "000000";
				when "000100000011" => data <= "000000";
				when "000100000100" => data <= "000000";
				when "000100000101" => data <= "000000";
				when "000100000110" => data <= "000000";
				when "000100000111" => data <= "000000";
				when "000100001000" => data <= "000000";
				when "000100001001" => data <= "000000";
				when "000100001010" => data <= "000000";
				when "000100001011" => data <= "000000";
				when "000100001100" => data <= "000000";
				when "000100001101" => data <= "000000";
				when "000100001110" => data <= "000000";
				when "000100001111" => data <= "000000";
				when "000100010000" => data <= "000000";
				when "000100010001" => data <= "000000";
				when "000100010010" => data <= "000000";
				when "000100010011" => data <= "000000";
				when "000100010100" => data <= "000000";
				when "000100010101" => data <= "000000";
				when "000100010110" => data <= "000000";
				when "000100010111" => data <= "000000";
				when "000100011000" => data <= "000000";
				when "000100011001" => data <= "000000";
				when "000100011010" => data <= "000000";
				when "000100011011" => data <= "000000";
				when "000100011100" => data <= "000000";
				when "000100011101" => data <= "000000";
				when "000100011110" => data <= "000000";
				when "000100011111" => data <= "000000";
				when "000100100000" => data <= "000000";
				when "000100100001" => data <= "000000";
				when "000100100010" => data <= "000000";
				when "000100100011" => data <= "000000";
				when "000100100100" => data <= "000000";
				when "000100100101" => data <= "000000";
				when "000100100110" => data <= "000000";
				when "000100100111" => data <= "000000";
				when "000100101000" => data <= "000000";
				when "000100101001" => data <= "000000";
				when "000100101010" => data <= "000000";
				when "000100101011" => data <= "000000";
				when "000100101100" => data <= "000000";
				when "000100101101" => data <= "000000";
				when "000100101110" => data <= "000000";
				when "000100101111" => data <= "000000";
				when "000100110000" => data <= "000000";
				when "000100110001" => data <= "000000";
				when "000100110010" => data <= "000000";
				when "000100110011" => data <= "000000";
				when "000100110100" => data <= "000000";
				when "000100110101" => data <= "000000";
				when "000100110110" => data <= "000000";
				when "000100110111" => data <= "000000";
				when "000100111000" => data <= "000000";
				when "000100111001" => data <= "000000";
				when "000100111010" => data <= "000000";
				when "000100111011" => data <= "000000";
				when "000100111100" => data <= "000000";
				when "000100111101" => data <= "000000";
				when "000100111110" => data <= "000000";
				when "000100111111" => data <= "000000";
				when "000101000000" => data <= "000000";
				when "000101000001" => data <= "000000";
				when "000101000010" => data <= "000000";
				when "000101000011" => data <= "000000";
				when "000101000100" => data <= "000000";
				when "000101000101" => data <= "000000";
				when "000101000110" => data <= "000000";
				when "000101000111" => data <= "000000";
				when "000101001000" => data <= "000000";
				when "000101001001" => data <= "000000";
				when "000101001010" => data <= "000000";
				when "000101001011" => data <= "000000";
				when "000101001100" => data <= "000000";
				when "000101001101" => data <= "000000";
				when "000101001110" => data <= "000000";
				when "000101001111" => data <= "000000";
				when "000101010000" => data <= "000000";
				when "000101010001" => data <= "000000";
				when "000101010010" => data <= "000000";
				when "000101010011" => data <= "000000";
				when "000101010100" => data <= "000000";
				when "000101010101" => data <= "000000";
				when "000101010110" => data <= "000000";
				when "000101010111" => data <= "000000";
				when "000101011000" => data <= "000000";
				when "000101011001" => data <= "000000";
				when "000101011010" => data <= "000000";
				when "000101011011" => data <= "000000";
				when "000101011100" => data <= "000000";
				when "000101011101" => data <= "000000";
				when "000101011110" => data <= "000000";
				when "000101011111" => data <= "000000";
				when "000101100000" => data <= "000000";
				when "000101100001" => data <= "000000";
				when "000101100010" => data <= "000000";
				when "000101100011" => data <= "000000";
				when "000101100100" => data <= "000000";
				when "000101100101" => data <= "000000";
				when "000101100110" => data <= "000000";
				when "000101100111" => data <= "000000";
				when "000101101000" => data <= "000000";
				when "000101101001" => data <= "000000";
				when "000101101010" => data <= "000000";
				when "000101101011" => data <= "000000";
				when "000101101100" => data <= "000000";
				when "000101101101" => data <= "000000";
				when "000101101110" => data <= "000000";
				when "000101101111" => data <= "000000";
				when "000101110000" => data <= "000000";
				when "000101110001" => data <= "000000";
				when "000101110010" => data <= "000000";
				when "000101110011" => data <= "000000";
				when "000101110100" => data <= "000000";
				when "000101110101" => data <= "000000";
				when "000101110110" => data <= "000000";
				when "000101110111" => data <= "000000";
				when "000101111000" => data <= "000000";
				when "000101111001" => data <= "000000";
				when "000101111010" => data <= "000000";
				when "000101111011" => data <= "000000";
				when "000101111100" => data <= "000000";
				when "000101111101" => data <= "000000";
				when "000101111110" => data <= "000000";
				when "000101111111" => data <= "000000";
				when "000110000000" => data <= "000000";
				when "000110000001" => data <= "000000";
				when "000110000010" => data <= "000000";
				when "000110000011" => data <= "000000";
				when "000110000100" => data <= "000000";
				when "000110000101" => data <= "000000";
				when "000110000110" => data <= "000000";
				when "000110000111" => data <= "000000";
				when "000110001000" => data <= "000000";
				when "000110001001" => data <= "000000";
				when "000110001010" => data <= "000000";
				when "000110001011" => data <= "000000";
				when "000110001100" => data <= "000000";
				when "000110001101" => data <= "000000";
				when "000110001110" => data <= "000000";
				when "000110001111" => data <= "000000";
				when "000110010000" => data <= "000000";
				when "000110010001" => data <= "000000";
				when "000110010010" => data <= "000000";
				when "000110010011" => data <= "000000";
				when "000110010100" => data <= "000000";
				when "000110010101" => data <= "000000";
				when "000110010110" => data <= "000000";
				when "000110010111" => data <= "000000";
				when "000110011000" => data <= "000000";
				when "000110011001" => data <= "000000";
				when "000110011010" => data <= "000000";
				when "000110011011" => data <= "000000";
				when "000110011100" => data <= "000000";
				when "000110011101" => data <= "000000";
				when "000110011110" => data <= "000000";
				when "000110011111" => data <= "000000";
				when "000110100000" => data <= "000000";
				when "000110100001" => data <= "000000";
				when "000110100010" => data <= "000000";
				when "000110100011" => data <= "000000";
				when "000110100100" => data <= "000000";
				when "000110100101" => data <= "000000";
				when "000110100110" => data <= "000000";
				when "000110100111" => data <= "000000";
				when "000110101000" => data <= "000000";
				when "000110101001" => data <= "000000";
				when "000110101010" => data <= "000000";
				when "000110101011" => data <= "000000";
				when "000110101100" => data <= "000000";
				when "000110101101" => data <= "000000";
				when "000110101110" => data <= "000000";
				when "000110101111" => data <= "000000";
				when "000110110000" => data <= "000000";
				when "000110110001" => data <= "000000";
				when "000110110010" => data <= "000000";
				when "000110110011" => data <= "000000";
				when "000110110100" => data <= "000000";
				when "000110110101" => data <= "000000";
				when "000110110110" => data <= "000000";
				when "000110110111" => data <= "000000";
				when "000110111000" => data <= "000000";
				when "000110111001" => data <= "000000";
				when "000110111010" => data <= "000000";
				when "000110111011" => data <= "000000";
				when "000110111100" => data <= "000000";
				when "000110111101" => data <= "000000";
				when "000110111110" => data <= "000000";
				when "000110111111" => data <= "000000";
				when "000111000000" => data <= "000000";
				when "000111000001" => data <= "000000";
				when "000111000010" => data <= "000000";
				when "000111000011" => data <= "000000";
				when "000111000100" => data <= "000000";
				when "000111000101" => data <= "000000";
				when "000111000110" => data <= "000000";
				when "000111000111" => data <= "000000";
				when "000111001000" => data <= "000000";
				when "000111001001" => data <= "000000";
				when "000111001010" => data <= "000000";
				when "000111001011" => data <= "000000";
				when "000111001100" => data <= "000000";
				when "000111001101" => data <= "000000";
				when "000111001110" => data <= "000000";
				when "000111001111" => data <= "000000";
				when "000111010000" => data <= "000000";
				when "000111010001" => data <= "000000";
				when "000111010010" => data <= "000000";
				when "000111010011" => data <= "000000";
				when "000111010100" => data <= "000000";
				when "000111010101" => data <= "000000";
				when "000111010110" => data <= "000000";
				when "000111010111" => data <= "000000";
				when "000111011000" => data <= "000000";
				when "000111011001" => data <= "000000";
				when "000111011010" => data <= "000000";
				when "000111011011" => data <= "000000";
				when "000111011100" => data <= "000000";
				when "000111011101" => data <= "000000";
				when "000111011110" => data <= "000000";
				when "000111011111" => data <= "000000";
				when "000111100000" => data <= "000000";
				when "000111100001" => data <= "000000";
				when "000111100010" => data <= "000000";
				when "000111100011" => data <= "000000";
				when "000111100100" => data <= "000000";
				when "000111100101" => data <= "000000";
				when "000111100110" => data <= "000000";
				when "000111100111" => data <= "000000";
				when "000111101000" => data <= "000000";
				when "000111101001" => data <= "000000";
				when "000111101010" => data <= "000000";
				when "000111101011" => data <= "000000";
				when "000111101100" => data <= "000000";
				when "000111101101" => data <= "000000";
				when "000111101110" => data <= "000000";
				when "000111101111" => data <= "000000";
				when "000111110000" => data <= "000000";
				when "000111110001" => data <= "000000";
				when "000111110010" => data <= "000000";
				when "000111110011" => data <= "000000";
				when "000111110100" => data <= "000000";
				when "000111110101" => data <= "000000";
				when "000111110110" => data <= "000000";
				when "000111110111" => data <= "000000";
				when "000111111000" => data <= "000000";
				when "000111111001" => data <= "000000";
				when "000111111010" => data <= "000000";
				when "000111111011" => data <= "000000";
				when "000111111100" => data <= "000000";
				when "000111111101" => data <= "000000";
				when "000111111110" => data <= "000000";
				when "000111111111" => data <= "000000";
				when "001000000000" => data <= "000000";
				when "001000000001" => data <= "000000";
				when "001000000010" => data <= "000000";
				when "001000000011" => data <= "000000";
				when "001000000100" => data <= "000000";
				when "001000000101" => data <= "000000";
				when "001000000110" => data <= "000000";
				when "001000000111" => data <= "000000";
				when "001000001000" => data <= "000000";
				when "001000001001" => data <= "000000";
				when "001000001010" => data <= "000000";
				when "001000001011" => data <= "000000";
				when "001000001100" => data <= "000000";
				when "001000001101" => data <= "000000";
				when "001000001110" => data <= "000000";
				when "001000001111" => data <= "000000";
				when "001000010000" => data <= "000000";
				when "001000010001" => data <= "000000";
				when "001000010010" => data <= "000000";
				when "001000010011" => data <= "000000";
				when "001000010100" => data <= "000000";
				when "001000010101" => data <= "000000";
				when "001000010110" => data <= "000000";
				when "001000010111" => data <= "000000";
				when "001000011000" => data <= "000000";
				when "001000011001" => data <= "000000";
				when "001000011010" => data <= "000000";
				when "001000011011" => data <= "000000";
				when "001000011100" => data <= "000000";
				when "001000011101" => data <= "000000";
				when "001000011110" => data <= "000000";
				when "001000011111" => data <= "000000";
				when "001000100000" => data <= "000000";
				when "001000100001" => data <= "000000";
				when "001000100010" => data <= "000000";
				when "001000100011" => data <= "000000";
				when "001000100100" => data <= "000000";
				when "001000100101" => data <= "000000";
				when "001000100110" => data <= "000000";
				when "001000100111" => data <= "000000";
				when "001000101000" => data <= "000000";
				when "001000101001" => data <= "000000";
				when "001000101010" => data <= "000000";
				when "001000101011" => data <= "000000";
				when "001000101100" => data <= "000000";
				when "001000101101" => data <= "000000";
				when "001000101110" => data <= "000000";
				when "001000101111" => data <= "000000";
				when "001000110000" => data <= "000000";
				when "001000110001" => data <= "000000";
				when "001000110010" => data <= "000000";
				when "001000110011" => data <= "000000";
				when "001000110100" => data <= "000000";
				when "001000110101" => data <= "000000";
				when "001000110110" => data <= "000000";
				when "001000110111" => data <= "000000";
				when "001000111000" => data <= "000000";
				when "001000111001" => data <= "000000";
				when "001000111010" => data <= "000000";
				when "001000111011" => data <= "000000";
				when "001000111100" => data <= "000000";
				when "001000111101" => data <= "000000";
				when "001000111110" => data <= "000000";
				when "001000111111" => data <= "000000";
				when "001001000000" => data <= "000000";
				when "001001000001" => data <= "000000";
				when "001001000010" => data <= "000000";
				when "001001000011" => data <= "000000";
				when "001001000100" => data <= "000000";
				when "001001000101" => data <= "000000";
				when "001001000110" => data <= "000000";
				when "001001000111" => data <= "000000";
				when "001001001000" => data <= "000000";
				when "001001001001" => data <= "000000";
				when "001001001010" => data <= "000000";
				when "001001001011" => data <= "000000";
				when "001001001100" => data <= "000000";
				when "001001001101" => data <= "000000";
				when "001001001110" => data <= "000000";
				when "001001001111" => data <= "000000";
				when "001001010000" => data <= "000000";
				when "001001010001" => data <= "000000";
				when "001001010010" => data <= "000000";
				when "001001010011" => data <= "000000";
				when "001001010100" => data <= "000000";
				when "001001010101" => data <= "000000";
				when "001001010110" => data <= "000000";
				when "001001010111" => data <= "000000";
				when "001001011000" => data <= "000000";
				when "001001011001" => data <= "000000";
				when "001001011010" => data <= "000000";
				when "001001011011" => data <= "000000";
				when "001001011100" => data <= "000000";
				when "001001011101" => data <= "000000";
				when "001001011110" => data <= "000000";
				when "001001011111" => data <= "000000";
				when "001001100000" => data <= "000000";
				when "001001100001" => data <= "000000";
				when "001001100010" => data <= "000000";
				when "001001100011" => data <= "000000";
				when "001001100100" => data <= "000000";
				when "001001100101" => data <= "000000";
				when "001001100110" => data <= "000000";
				when "001001100111" => data <= "000000";
				when "001001101000" => data <= "000000";
				when "001001101001" => data <= "000000";
				when "001001101010" => data <= "000000";
				when "001001101011" => data <= "000000";
				when "001001101100" => data <= "000000";
				when "001001101101" => data <= "000000";
				when "001001101110" => data <= "000000";
				when "001001101111" => data <= "000000";
				when "001001110000" => data <= "000000";
				when "001001110001" => data <= "000000";
				when "001001110010" => data <= "000000";
				when "001001110011" => data <= "000000";
				when "001001110100" => data <= "000000";
				when "001001110101" => data <= "000000";
				when "001001110110" => data <= "000000";
				when "001001110111" => data <= "000000";
				when "001001111000" => data <= "000000";
				when "001001111001" => data <= "000000";
				when "001001111010" => data <= "000000";
				when "001001111011" => data <= "000000";
				when "001001111100" => data <= "000000";
				when "001001111101" => data <= "000000";
				when "001001111110" => data <= "000000";
				when "001001111111" => data <= "000000";
				when "001010000000" => data <= "000000";
				when "001010000001" => data <= "000000";
				when "001010000010" => data <= "000000";
				when "001010000011" => data <= "000000";
				when "001010000100" => data <= "000000";
				when "001010000101" => data <= "000000";
				when "001010000110" => data <= "000000";
				when "001010000111" => data <= "000000";
				when "001010001000" => data <= "000000";
				when "001010001001" => data <= "000000";
				when "001010001010" => data <= "000000";
				when "001010001011" => data <= "000000";
				when "001010001100" => data <= "000000";
				when "001010001101" => data <= "000000";
				when "001010001110" => data <= "000000";
				when "001010001111" => data <= "000000";
				when "001010010000" => data <= "000000";
				when "001010010001" => data <= "000000";
				when "001010010010" => data <= "000000";
				when "001010010011" => data <= "000000";
				when "001010010100" => data <= "000000";
				when "001010010101" => data <= "000000";
				when "001010010110" => data <= "000000";
				when "001010010111" => data <= "000000";
				when "001010011000" => data <= "000000";
				when "001010011001" => data <= "000000";
				when "001010011010" => data <= "000000";
				when "001010011011" => data <= "000000";
				when "001010011100" => data <= "000000";
				when "001010011101" => data <= "000000";
				when "001010011110" => data <= "000000";
				when "001010011111" => data <= "000000";
				when "001010100000" => data <= "000000";
				when "001010100001" => data <= "000000";
				when "001010100010" => data <= "000000";
				when "001010100011" => data <= "000000";
				when "001010100100" => data <= "000000";
				when "001010100101" => data <= "000000";
				when "001010100110" => data <= "000000";
				when "001010100111" => data <= "000000";
				when "001010101000" => data <= "000000";
				when "001010101001" => data <= "000000";
				when "001010101010" => data <= "000000";
				when "001010101011" => data <= "000000";
				when "001010101100" => data <= "000000";
				when "001010101101" => data <= "000000";
				when "001010101110" => data <= "000000";
				when "001010101111" => data <= "000000";
				when "001010110000" => data <= "000000";
				when "001010110001" => data <= "000000";
				when "001010110010" => data <= "000000";
				when "001010110011" => data <= "000000";
				when "001010110100" => data <= "000000";
				when "001010110101" => data <= "000000";
				when "001010110110" => data <= "000000";
				when "001010110111" => data <= "000000";
				when "001010111000" => data <= "000000";
				when "001010111001" => data <= "000000";
				when "001010111010" => data <= "000000";
				when "001010111011" => data <= "000000";
				when "001010111100" => data <= "000000";
				when "001010111101" => data <= "000000";
				when "001010111110" => data <= "000000";
				when "001010111111" => data <= "000000";
				when "001011000000" => data <= "000000";
				when "001011000001" => data <= "000000";
				when "001011000010" => data <= "000000";
				when "001011000011" => data <= "000000";
				when "001011000100" => data <= "000000";
				when "001011000101" => data <= "000000";
				when "001011000110" => data <= "000000";
				when "001011000111" => data <= "000000";
				when "001011001000" => data <= "000000";
				when "001011001001" => data <= "000000";
				when "001011001010" => data <= "000000";
				when "001011001011" => data <= "000000";
				when "001011001100" => data <= "000000";
				when "001011001101" => data <= "000000";
				when "001011001110" => data <= "000000";
				when "001011001111" => data <= "000000";
				when "001011010000" => data <= "000000";
				when "001011010001" => data <= "000000";
				when "001011010010" => data <= "000000";
				when "001011010011" => data <= "000000";
				when "001011010100" => data <= "000000";
				when "001011010101" => data <= "000000";
				when "001011010110" => data <= "000000";
				when "001011010111" => data <= "000000";
				when "001011011000" => data <= "000000";
				when "001011011001" => data <= "000000";
				when "001011011010" => data <= "000000";
				when "001011011011" => data <= "000000";
				when "001011011100" => data <= "000000";
				when "001011011101" => data <= "000000";
				when "001011011110" => data <= "000000";
				when "001011011111" => data <= "000000";
				when "001011100000" => data <= "000000";
				when "001011100001" => data <= "000000";
				when "001011100010" => data <= "000000";
				when "001011100011" => data <= "000000";
				when "001011100100" => data <= "000000";
				when "001011100101" => data <= "000000";
				when "001011100110" => data <= "000000";
				when "001011100111" => data <= "000000";
				when "001011101000" => data <= "000000";
				when "001011101001" => data <= "000000";
				when "001011101010" => data <= "000000";
				when "001011101011" => data <= "000000";
				when "001011101100" => data <= "000000";
				when "001011101101" => data <= "000000";
				when "001011101110" => data <= "000000";
				when "001011101111" => data <= "000000";
				when "001011110000" => data <= "000000";
				when "001011110001" => data <= "000000";
				when "001011110010" => data <= "000000";
				when "001011110011" => data <= "000000";
				when "001011110100" => data <= "000000";
				when "001011110101" => data <= "000000";
				when "001011110110" => data <= "000000";
				when "001011110111" => data <= "000000";
				when "001011111000" => data <= "000000";
				when "001011111001" => data <= "000000";
				when "001011111010" => data <= "000000";
				when "001011111011" => data <= "000000";
				when "001011111100" => data <= "000000";
				when "001011111101" => data <= "000000";
				when "001011111110" => data <= "000000";
				when "001011111111" => data <= "000000";
				when "001100000000" => data <= "000000";
				when "001100000001" => data <= "000000";
				when "001100000010" => data <= "000000";
				when "001100000011" => data <= "000000";
				when "001100000100" => data <= "000000";
				when "001100000101" => data <= "000000";
				when "001100000110" => data <= "000000";
				when "001100000111" => data <= "000000";
				when "001100001000" => data <= "000000";
				when "001100001001" => data <= "000000";
				when "001100001010" => data <= "000000";
				when "001100001011" => data <= "000000";
				when "001100001100" => data <= "000000";
				when "001100001101" => data <= "000000";
				when "001100001110" => data <= "000000";
				when "001100001111" => data <= "000000";
				when "001100010000" => data <= "000000";
				when "001100010001" => data <= "000000";
				when "001100010010" => data <= "000000";
				when "001100010011" => data <= "000000";
				when "001100010100" => data <= "000000";
				when "001100010101" => data <= "111111";
				when "001100010110" => data <= "111111";
				when "001100010111" => data <= "111111";
				when "001100011000" => data <= "111111";
				when "001100011001" => data <= "111111";
				when "001100011010" => data <= "111111";
				when "001100011011" => data <= "111111";
				when "001100011100" => data <= "111111";
				when "001100011101" => data <= "000000";
				when "001100011110" => data <= "000000";
				when "001100011111" => data <= "000000";
				when "001100100000" => data <= "000000";
				when "001100100001" => data <= "000000";
				when "001100100010" => data <= "000000";
				when "001100100011" => data <= "000000";
				when "001100100100" => data <= "000000";
				when "001100100101" => data <= "000000";
				when "001100100110" => data <= "000000";
				when "001100100111" => data <= "111111";
				when "001100101000" => data <= "111111";
				when "001100101001" => data <= "111111";
				when "001100101010" => data <= "111111";
				when "001100101011" => data <= "111111";
				when "001100101100" => data <= "111111";
				when "001100101101" => data <= "111111";
				when "001100101110" => data <= "111111";
				when "001100101111" => data <= "111111";
				when "001100110000" => data <= "111111";
				when "001100110001" => data <= "000000";
				when "001100110010" => data <= "000000";
				when "001100110011" => data <= "000000";
				when "001100110100" => data <= "000000";
				when "001100110101" => data <= "000000";
				when "001100110110" => data <= "000000";
				when "001100110111" => data <= "000000";
				when "001100111000" => data <= "111111";
				when "001100111001" => data <= "111111";
				when "001100111010" => data <= "111111";
				when "001100111011" => data <= "111111";
				when "001100111100" => data <= "111111";
				when "001100111101" => data <= "111111";
				when "001100111110" => data <= "111111";
				when "001100111111" => data <= "111111";
				when "001101000000" => data <= "111111";
				when "001101000001" => data <= "111111";
				when "001101000010" => data <= "111111";
				when "001101000011" => data <= "111111";
				when "001101000100" => data <= "000000";
				when "001101000101" => data <= "000000";
				when "001101000110" => data <= "000000";
				when "001101000111" => data <= "000000";
				when "001101001000" => data <= "000000";
				when "001101001001" => data <= "000000";
				when "001101001010" => data <= "000000";
				when "001101001011" => data <= "111111";
				when "001101001100" => data <= "111111";
				when "001101001101" => data <= "111111";
				when "001101001110" => data <= "111111";
				when "001101001111" => data <= "111111";
				when "001101010000" => data <= "111111";
				when "001101010001" => data <= "111111";
				when "001101010010" => data <= "111111";
				when "001101010011" => data <= "000000";
				when "001101010100" => data <= "000000";
				when "001101010101" => data <= "000000";
				when "001101010110" => data <= "000000";
				when "001101010111" => data <= "000000";
				when "001101011000" => data <= "000000";
				when "001101011001" => data <= "000000";
				when "001101011010" => data <= "000000";
				when "001101011011" => data <= "000000";
				when "001101011100" => data <= "000000";
				when "001101011101" => data <= "000000";
				when "001101011110" => data <= "111111";
				when "001101011111" => data <= "111111";
				when "001101100000" => data <= "111111";
				when "001101100001" => data <= "111111";
				when "001101100010" => data <= "111111";
				when "001101100011" => data <= "111111";
				when "001101100100" => data <= "111111";
				when "001101100101" => data <= "111111";
				when "001101100110" => data <= "000000";
				when "001101100111" => data <= "000000";
				when "001101101000" => data <= "000000";
				when "001101101001" => data <= "000000";
				when "001101101010" => data <= "000000";
				when "001101101011" => data <= "000000";
				when "001101101100" => data <= "000000";
				when "001101101101" => data <= "000000";
				when "001101101110" => data <= "000000";
				when "001101101111" => data <= "000000";
				when "001101110000" => data <= "000000";
				when "001101110001" => data <= "000000";
				when "001101110010" => data <= "000000";
				when "001101110011" => data <= "000000";
				when "001101110100" => data <= "000000";
				when "001101110101" => data <= "000000";
				when "001101110110" => data <= "000000";
				when "001101110111" => data <= "000000";
				when "001101111000" => data <= "000000";
				when "001101111001" => data <= "000000";
				when "001101111010" => data <= "000000";
				when "001101111011" => data <= "000000";
				when "001101111100" => data <= "000000";
				when "001101111101" => data <= "000000";
				when "001101111110" => data <= "000000";
				when "001101111111" => data <= "000000";
				when "001110000000" => data <= "000000";
				when "001110000001" => data <= "000000";
				when "001110000010" => data <= "000000";
				when "001110000011" => data <= "000000";
				when "001110000100" => data <= "000000";
				when "001110000101" => data <= "000000";
				when "001110000110" => data <= "000000";
				when "001110000111" => data <= "000000";
				when "001110001000" => data <= "000000";
				when "001110001001" => data <= "000000";
				when "001110001010" => data <= "000000";
				when "001110001011" => data <= "000000";
				when "001110001100" => data <= "000000";
				when "001110001101" => data <= "000000";
				when "001110001110" => data <= "000000";
				when "001110001111" => data <= "000000";
				when "001110010000" => data <= "000000";
				when "001110010001" => data <= "000000";
				when "001110010010" => data <= "000000";
				when "001110010011" => data <= "000000";
				when "001110010100" => data <= "111111";
				when "001110010101" => data <= "010010";
				when "001110010110" => data <= "010010";
				when "001110010111" => data <= "010010";
				when "001110011000" => data <= "010010";
				when "001110011001" => data <= "010010";
				when "001110011010" => data <= "010010";
				when "001110011011" => data <= "010010";
				when "001110011100" => data <= "010010";
				when "001110011101" => data <= "111111";
				when "001110011110" => data <= "000000";
				when "001110011111" => data <= "000000";
				when "001110100000" => data <= "000000";
				when "001110100001" => data <= "000000";
				when "001110100010" => data <= "000000";
				when "001110100011" => data <= "000000";
				when "001110100100" => data <= "000000";
				when "001110100101" => data <= "000000";
				when "001110100110" => data <= "111111";
				when "001110100111" => data <= "010010";
				when "001110101000" => data <= "010010";
				when "001110101001" => data <= "010010";
				when "001110101010" => data <= "010010";
				when "001110101011" => data <= "010010";
				when "001110101100" => data <= "010010";
				when "001110101101" => data <= "010010";
				when "001110101110" => data <= "010010";
				when "001110101111" => data <= "010010";
				when "001110110000" => data <= "010010";
				when "001110110001" => data <= "111111";
				when "001110110010" => data <= "000000";
				when "001110110011" => data <= "000000";
				when "001110110100" => data <= "000000";
				when "001110110101" => data <= "000000";
				when "001110110110" => data <= "000000";
				when "001110110111" => data <= "111111";
				when "001110111000" => data <= "010010";
				when "001110111001" => data <= "010010";
				when "001110111010" => data <= "010010";
				when "001110111011" => data <= "010010";
				when "001110111100" => data <= "010010";
				when "001110111101" => data <= "010010";
				when "001110111110" => data <= "010010";
				when "001110111111" => data <= "010010";
				when "001111000000" => data <= "010010";
				when "001111000001" => data <= "010010";
				when "001111000010" => data <= "010010";
				when "001111000011" => data <= "010010";
				when "001111000100" => data <= "111111";
				when "001111000101" => data <= "000000";
				when "001111000110" => data <= "000000";
				when "001111000111" => data <= "000000";
				when "001111001000" => data <= "000000";
				when "001111001001" => data <= "000000";
				when "001111001010" => data <= "111111";
				when "001111001011" => data <= "010010";
				when "001111001100" => data <= "010010";
				when "001111001101" => data <= "010010";
				when "001111001110" => data <= "010010";
				when "001111001111" => data <= "010010";
				when "001111010000" => data <= "010010";
				when "001111010001" => data <= "010010";
				when "001111010010" => data <= "010010";
				when "001111010011" => data <= "111111";
				when "001111010100" => data <= "000000";
				when "001111010101" => data <= "000000";
				when "001111010110" => data <= "000000";
				when "001111010111" => data <= "000000";
				when "001111011000" => data <= "000000";
				when "001111011001" => data <= "000000";
				when "001111011010" => data <= "000000";
				when "001111011011" => data <= "000000";
				when "001111011100" => data <= "000000";
				when "001111011101" => data <= "111111";
				when "001111011110" => data <= "010010";
				when "001111011111" => data <= "010010";
				when "001111100000" => data <= "010010";
				when "001111100001" => data <= "010010";
				when "001111100010" => data <= "010010";
				when "001111100011" => data <= "010010";
				when "001111100100" => data <= "010010";
				when "001111100101" => data <= "010010";
				when "001111100110" => data <= "111111";
				when "001111100111" => data <= "000000";
				when "001111101000" => data <= "000000";
				when "001111101001" => data <= "000000";
				when "001111101010" => data <= "000000";
				when "001111101011" => data <= "000000";
				when "001111101100" => data <= "000000";
				when "001111101101" => data <= "000000";
				when "001111101110" => data <= "000000";
				when "001111101111" => data <= "000000";
				when "001111110000" => data <= "000000";
				when "001111110001" => data <= "000000";
				when "001111110010" => data <= "000000";
				when "001111110011" => data <= "000000";
				when "001111110100" => data <= "000000";
				when "001111110101" => data <= "000000";
				when "001111110110" => data <= "000000";
				when "001111110111" => data <= "000000";
				when "001111111000" => data <= "000000";
				when "001111111001" => data <= "000000";
				when "001111111010" => data <= "000000";
				when "001111111011" => data <= "000000";
				when "001111111100" => data <= "000000";
				when "001111111101" => data <= "000000";
				when "001111111110" => data <= "000000";
				when "001111111111" => data <= "000000";
				when "010000000000" => data <= "000000";
				when "010000000001" => data <= "000000";
				when "010000000010" => data <= "000000";
				when "010000000011" => data <= "000000";
				when "010000000100" => data <= "000000";
				when "010000000101" => data <= "000000";
				when "010000000110" => data <= "000000";
				when "010000000111" => data <= "000000";
				when "010000001000" => data <= "000000";
				when "010000001001" => data <= "000000";
				when "010000001010" => data <= "000000";
				when "010000001011" => data <= "000000";
				when "010000001100" => data <= "000000";
				when "010000001101" => data <= "000000";
				when "010000001110" => data <= "000000";
				when "010000001111" => data <= "000000";
				when "010000010000" => data <= "000000";
				when "010000010001" => data <= "000000";
				when "010000010010" => data <= "000000";
				when "010000010011" => data <= "000000";
				when "010000010100" => data <= "111111";
				when "010000010101" => data <= "010010";
				when "010000010110" => data <= "010010";
				when "010000010111" => data <= "010010";
				when "010000011000" => data <= "010010";
				when "010000011001" => data <= "010010";
				when "010000011010" => data <= "010010";
				when "010000011011" => data <= "010010";
				when "010000011100" => data <= "010010";
				when "010000011101" => data <= "111111";
				when "010000011110" => data <= "111111";
				when "010000011111" => data <= "000000";
				when "010000100000" => data <= "000000";
				when "010000100001" => data <= "000000";
				when "010000100010" => data <= "000000";
				when "010000100011" => data <= "000000";
				when "010000100100" => data <= "000000";
				when "010000100101" => data <= "000000";
				when "010000100110" => data <= "111111";
				when "010000100111" => data <= "010010";
				when "010000101000" => data <= "010010";
				when "010000101001" => data <= "010010";
				when "010000101010" => data <= "010010";
				when "010000101011" => data <= "010010";
				when "010000101100" => data <= "010010";
				when "010000101101" => data <= "010010";
				when "010000101110" => data <= "010010";
				when "010000101111" => data <= "010010";
				when "010000110000" => data <= "010010";
				when "010000110001" => data <= "111111";
				when "010000110010" => data <= "000000";
				when "010000110011" => data <= "000000";
				when "010000110100" => data <= "000000";
				when "010000110101" => data <= "000000";
				when "010000110110" => data <= "000000";
				when "010000110111" => data <= "111111";
				when "010000111000" => data <= "010010";
				when "010000111001" => data <= "010010";
				when "010000111010" => data <= "010010";
				when "010000111011" => data <= "010010";
				when "010000111100" => data <= "010010";
				when "010000111101" => data <= "010010";
				when "010000111110" => data <= "010010";
				when "010000111111" => data <= "010010";
				when "010001000000" => data <= "010010";
				when "010001000001" => data <= "010010";
				when "010001000010" => data <= "010010";
				when "010001000011" => data <= "010010";
				when "010001000100" => data <= "111111";
				when "010001000101" => data <= "000000";
				when "010001000110" => data <= "000000";
				when "010001000111" => data <= "000000";
				when "010001001000" => data <= "000000";
				when "010001001001" => data <= "000000";
				when "010001001010" => data <= "111111";
				when "010001001011" => data <= "010010";
				when "010001001100" => data <= "010010";
				when "010001001101" => data <= "010010";
				when "010001001110" => data <= "010010";
				when "010001001111" => data <= "010010";
				when "010001010000" => data <= "010010";
				when "010001010001" => data <= "010010";
				when "010001010010" => data <= "010010";
				when "010001010011" => data <= "111111";
				when "010001010100" => data <= "111111";
				when "010001010101" => data <= "000000";
				when "010001010110" => data <= "000000";
				when "010001010111" => data <= "000000";
				when "010001011000" => data <= "000000";
				when "010001011001" => data <= "000000";
				when "010001011010" => data <= "000000";
				when "010001011011" => data <= "000000";
				when "010001011100" => data <= "111111";
				when "010001011101" => data <= "010010";
				when "010001011110" => data <= "010010";
				when "010001011111" => data <= "010010";
				when "010001100000" => data <= "010010";
				when "010001100001" => data <= "010010";
				when "010001100010" => data <= "010010";
				when "010001100011" => data <= "010010";
				when "010001100100" => data <= "010010";
				when "010001100101" => data <= "010010";
				when "010001100110" => data <= "010010";
				when "010001100111" => data <= "111111";
				when "010001101000" => data <= "000000";
				when "010001101001" => data <= "000000";
				when "010001101010" => data <= "000000";
				when "010001101011" => data <= "000000";
				when "010001101100" => data <= "000000";
				when "010001101101" => data <= "000000";
				when "010001101110" => data <= "000000";
				when "010001101111" => data <= "000000";
				when "010001110000" => data <= "000000";
				when "010001110001" => data <= "000000";
				when "010001110010" => data <= "000000";
				when "010001110011" => data <= "000000";
				when "010001110100" => data <= "000000";
				when "010001110101" => data <= "000000";
				when "010001110110" => data <= "000000";
				when "010001110111" => data <= "000000";
				when "010001111000" => data <= "000000";
				when "010001111001" => data <= "000000";
				when "010001111010" => data <= "000000";
				when "010001111011" => data <= "000000";
				when "010001111100" => data <= "000000";
				when "010001111101" => data <= "000000";
				when "010001111110" => data <= "000000";
				when "010001111111" => data <= "000000";
				when "010010000000" => data <= "000000";
				when "010010000001" => data <= "000000";
				when "010010000010" => data <= "000000";
				when "010010000011" => data <= "000000";
				when "010010000100" => data <= "000000";
				when "010010000101" => data <= "000000";
				when "010010000110" => data <= "000000";
				when "010010000111" => data <= "000000";
				when "010010001000" => data <= "000000";
				when "010010001001" => data <= "000000";
				when "010010001010" => data <= "000000";
				when "010010001011" => data <= "000000";
				when "010010001100" => data <= "000000";
				when "010010001101" => data <= "000000";
				when "010010001110" => data <= "000000";
				when "010010001111" => data <= "000000";
				when "010010010000" => data <= "000000";
				when "010010010001" => data <= "000000";
				when "010010010010" => data <= "000000";
				when "010010010011" => data <= "000000";
				when "010010010100" => data <= "111111";
				when "010010010101" => data <= "010010";
				when "010010010110" => data <= "010010";
				when "010010010111" => data <= "111111";
				when "010010011000" => data <= "111111";
				when "010010011001" => data <= "111111";
				when "010010011010" => data <= "111111";
				when "010010011011" => data <= "111111";
				when "010010011100" => data <= "111111";
				when "010010011101" => data <= "010010";
				when "010010011110" => data <= "010010";
				when "010010011111" => data <= "111111";
				when "010010100000" => data <= "000000";
				when "010010100001" => data <= "000000";
				when "010010100010" => data <= "000000";
				when "010010100011" => data <= "000000";
				when "010010100100" => data <= "000000";
				when "010010100101" => data <= "000000";
				when "010010100110" => data <= "111111";
				when "010010100111" => data <= "010010";
				when "010010101000" => data <= "010010";
				when "010010101001" => data <= "111111";
				when "010010101010" => data <= "111111";
				when "010010101011" => data <= "111111";
				when "010010101100" => data <= "111111";
				when "010010101101" => data <= "111111";
				when "010010101110" => data <= "111111";
				when "010010101111" => data <= "111111";
				when "010010110000" => data <= "111111";
				when "010010110001" => data <= "000000";
				when "010010110010" => data <= "000000";
				when "010010110011" => data <= "000000";
				when "010010110100" => data <= "000000";
				when "010010110101" => data <= "000000";
				when "010010110110" => data <= "000000";
				when "010010110111" => data <= "000000";
				when "010010111000" => data <= "111111";
				when "010010111001" => data <= "111111";
				when "010010111010" => data <= "111111";
				when "010010111011" => data <= "111111";
				when "010010111100" => data <= "111111";
				when "010010111101" => data <= "010010";
				when "010010111110" => data <= "010010";
				when "010010111111" => data <= "111111";
				when "010011000000" => data <= "111111";
				when "010011000001" => data <= "111111";
				when "010011000010" => data <= "111111";
				when "010011000011" => data <= "111111";
				when "010011000100" => data <= "000000";
				when "010011000101" => data <= "000000";
				when "010011000110" => data <= "000000";
				when "010011000111" => data <= "000000";
				when "010011001000" => data <= "000000";
				when "010011001001" => data <= "000000";
				when "010011001010" => data <= "111111";
				when "010011001011" => data <= "010010";
				when "010011001100" => data <= "010010";
				when "010011001101" => data <= "111111";
				when "010011001110" => data <= "111111";
				when "010011001111" => data <= "111111";
				when "010011010000" => data <= "111111";
				when "010011010001" => data <= "111111";
				when "010011010010" => data <= "111111";
				when "010011010011" => data <= "010010";
				when "010011010100" => data <= "010010";
				when "010011010101" => data <= "111111";
				when "010011010110" => data <= "000000";
				when "010011010111" => data <= "000000";
				when "010011011000" => data <= "000000";
				when "010011011001" => data <= "000000";
				when "010011011010" => data <= "000000";
				when "010011011011" => data <= "111111";
				when "010011011100" => data <= "010010";
				when "010011011101" => data <= "010010";
				when "010011011110" => data <= "111111";
				when "010011011111" => data <= "111111";
				when "010011100000" => data <= "111111";
				when "010011100001" => data <= "111111";
				when "010011100010" => data <= "111111";
				when "010011100011" => data <= "111111";
				when "010011100100" => data <= "111111";
				when "010011100101" => data <= "111111";
				when "010011100110" => data <= "010010";
				when "010011100111" => data <= "010010";
				when "010011101000" => data <= "111111";
				when "010011101001" => data <= "000000";
				when "010011101010" => data <= "000000";
				when "010011101011" => data <= "000000";
				when "010011101100" => data <= "000000";
				when "010011101101" => data <= "000000";
				when "010011101110" => data <= "000000";
				when "010011101111" => data <= "000000";
				when "010011110000" => data <= "000000";
				when "010011110001" => data <= "000000";
				when "010011110010" => data <= "000000";
				when "010011110011" => data <= "000000";
				when "010011110100" => data <= "000000";
				when "010011110101" => data <= "000000";
				when "010011110110" => data <= "000000";
				when "010011110111" => data <= "000000";
				when "010011111000" => data <= "000000";
				when "010011111001" => data <= "000000";
				when "010011111010" => data <= "000000";
				when "010011111011" => data <= "000000";
				when "010011111100" => data <= "000000";
				when "010011111101" => data <= "000000";
				when "010011111110" => data <= "000000";
				when "010011111111" => data <= "000000";
				when "010100000000" => data <= "000000";
				when "010100000001" => data <= "000000";
				when "010100000010" => data <= "000000";
				when "010100000011" => data <= "000000";
				when "010100000100" => data <= "000000";
				when "010100000101" => data <= "000000";
				when "010100000110" => data <= "000000";
				when "010100000111" => data <= "000000";
				when "010100001000" => data <= "000000";
				when "010100001001" => data <= "000000";
				when "010100001010" => data <= "000000";
				when "010100001011" => data <= "000000";
				when "010100001100" => data <= "000000";
				when "010100001101" => data <= "000000";
				when "010100001110" => data <= "000000";
				when "010100001111" => data <= "000000";
				when "010100010000" => data <= "000000";
				when "010100010001" => data <= "000000";
				when "010100010010" => data <= "000000";
				when "010100010011" => data <= "000000";
				when "010100010100" => data <= "111111";
				when "010100010101" => data <= "010010";
				when "010100010110" => data <= "010010";
				when "010100010111" => data <= "111111";
				when "010100011000" => data <= "000000";
				when "010100011001" => data <= "000000";
				when "010100011010" => data <= "000000";
				when "010100011011" => data <= "000000";
				when "010100011100" => data <= "111111";
				when "010100011101" => data <= "010010";
				when "010100011110" => data <= "010010";
				when "010100011111" => data <= "111111";
				when "010100100000" => data <= "000000";
				when "010100100001" => data <= "000000";
				when "010100100010" => data <= "000000";
				when "010100100011" => data <= "000000";
				when "010100100100" => data <= "000000";
				when "010100100101" => data <= "000000";
				when "010100100110" => data <= "111111";
				when "010100100111" => data <= "010010";
				when "010100101000" => data <= "010010";
				when "010100101001" => data <= "111111";
				when "010100101010" => data <= "000000";
				when "010100101011" => data <= "000000";
				when "010100101100" => data <= "000000";
				when "010100101101" => data <= "000000";
				when "010100101110" => data <= "000000";
				when "010100101111" => data <= "000000";
				when "010100110000" => data <= "000000";
				when "010100110001" => data <= "000000";
				when "010100110010" => data <= "000000";
				when "010100110011" => data <= "000000";
				when "010100110100" => data <= "000000";
				when "010100110101" => data <= "000000";
				when "010100110110" => data <= "000000";
				when "010100110111" => data <= "000000";
				when "010100111000" => data <= "000000";
				when "010100111001" => data <= "000000";
				when "010100111010" => data <= "000000";
				when "010100111011" => data <= "000000";
				when "010100111100" => data <= "111111";
				when "010100111101" => data <= "010010";
				when "010100111110" => data <= "010010";
				when "010100111111" => data <= "111111";
				when "010101000000" => data <= "000000";
				when "010101000001" => data <= "000000";
				when "010101000010" => data <= "000000";
				when "010101000011" => data <= "000000";
				when "010101000100" => data <= "000000";
				when "010101000101" => data <= "000000";
				when "010101000110" => data <= "000000";
				when "010101000111" => data <= "000000";
				when "010101001000" => data <= "000000";
				when "010101001001" => data <= "000000";
				when "010101001010" => data <= "111111";
				when "010101001011" => data <= "010010";
				when "010101001100" => data <= "010010";
				when "010101001101" => data <= "111111";
				when "010101001110" => data <= "000000";
				when "010101001111" => data <= "000000";
				when "010101010000" => data <= "000000";
				when "010101010001" => data <= "000000";
				when "010101010010" => data <= "111111";
				when "010101010011" => data <= "010010";
				when "010101010100" => data <= "010010";
				when "010101010101" => data <= "111111";
				when "010101010110" => data <= "000000";
				when "010101010111" => data <= "000000";
				when "010101011000" => data <= "000000";
				when "010101011001" => data <= "000000";
				when "010101011010" => data <= "000000";
				when "010101011011" => data <= "111111";
				when "010101011100" => data <= "010010";
				when "010101011101" => data <= "010010";
				when "010101011110" => data <= "111111";
				when "010101011111" => data <= "000000";
				when "010101100000" => data <= "000000";
				when "010101100001" => data <= "000000";
				when "010101100010" => data <= "000000";
				when "010101100011" => data <= "000000";
				when "010101100100" => data <= "000000";
				when "010101100101" => data <= "111111";
				when "010101100110" => data <= "010010";
				when "010101100111" => data <= "010010";
				when "010101101000" => data <= "111111";
				when "010101101001" => data <= "000000";
				when "010101101010" => data <= "000000";
				when "010101101011" => data <= "000000";
				when "010101101100" => data <= "000000";
				when "010101101101" => data <= "000000";
				when "010101101110" => data <= "000000";
				when "010101101111" => data <= "000000";
				when "010101110000" => data <= "000000";
				when "010101110001" => data <= "000000";
				when "010101110010" => data <= "000000";
				when "010101110011" => data <= "000000";
				when "010101110100" => data <= "000000";
				when "010101110101" => data <= "000000";
				when "010101110110" => data <= "000000";
				when "010101110111" => data <= "000000";
				when "010101111000" => data <= "000000";
				when "010101111001" => data <= "000000";
				when "010101111010" => data <= "000000";
				when "010101111011" => data <= "000000";
				when "010101111100" => data <= "000000";
				when "010101111101" => data <= "000000";
				when "010101111110" => data <= "000000";
				when "010101111111" => data <= "000000";
				when "010110000000" => data <= "000000";
				when "010110000001" => data <= "000000";
				when "010110000010" => data <= "000000";
				when "010110000011" => data <= "000000";
				when "010110000100" => data <= "000000";
				when "010110000101" => data <= "000000";
				when "010110000110" => data <= "000000";
				when "010110000111" => data <= "000000";
				when "010110001000" => data <= "000000";
				when "010110001001" => data <= "000000";
				when "010110001010" => data <= "000000";
				when "010110001011" => data <= "000000";
				when "010110001100" => data <= "000000";
				when "010110001101" => data <= "000000";
				when "010110001110" => data <= "000000";
				when "010110001111" => data <= "000000";
				when "010110010000" => data <= "000000";
				when "010110010001" => data <= "000000";
				when "010110010010" => data <= "000000";
				when "010110010011" => data <= "000000";
				when "010110010100" => data <= "111111";
				when "010110010101" => data <= "010010";
				when "010110010110" => data <= "010010";
				when "010110010111" => data <= "111111";
				when "010110011000" => data <= "000000";
				when "010110011001" => data <= "000000";
				when "010110011010" => data <= "000000";
				when "010110011011" => data <= "000000";
				when "010110011100" => data <= "111111";
				when "010110011101" => data <= "010010";
				when "010110011110" => data <= "010010";
				when "010110011111" => data <= "111111";
				when "010110100000" => data <= "000000";
				when "010110100001" => data <= "000000";
				when "010110100010" => data <= "000000";
				when "010110100011" => data <= "000000";
				when "010110100100" => data <= "000000";
				when "010110100101" => data <= "000000";
				when "010110100110" => data <= "111111";
				when "010110100111" => data <= "010010";
				when "010110101000" => data <= "010010";
				when "010110101001" => data <= "111111";
				when "010110101010" => data <= "000000";
				when "010110101011" => data <= "000000";
				when "010110101100" => data <= "000000";
				when "010110101101" => data <= "000000";
				when "010110101110" => data <= "000000";
				when "010110101111" => data <= "000000";
				when "010110110000" => data <= "000000";
				when "010110110001" => data <= "000000";
				when "010110110010" => data <= "000000";
				when "010110110011" => data <= "000000";
				when "010110110100" => data <= "000000";
				when "010110110101" => data <= "000000";
				when "010110110110" => data <= "000000";
				when "010110110111" => data <= "000000";
				when "010110111000" => data <= "000000";
				when "010110111001" => data <= "000000";
				when "010110111010" => data <= "000000";
				when "010110111011" => data <= "000000";
				when "010110111100" => data <= "111111";
				when "010110111101" => data <= "010010";
				when "010110111110" => data <= "010010";
				when "010110111111" => data <= "111111";
				when "010111000000" => data <= "000000";
				when "010111000001" => data <= "000000";
				when "010111000010" => data <= "000000";
				when "010111000011" => data <= "000000";
				when "010111000100" => data <= "000000";
				when "010111000101" => data <= "000000";
				when "010111000110" => data <= "000000";
				when "010111000111" => data <= "000000";
				when "010111001000" => data <= "000000";
				when "010111001001" => data <= "000000";
				when "010111001010" => data <= "111111";
				when "010111001011" => data <= "010010";
				when "010111001100" => data <= "010010";
				when "010111001101" => data <= "111111";
				when "010111001110" => data <= "000000";
				when "010111001111" => data <= "000000";
				when "010111010000" => data <= "000000";
				when "010111010001" => data <= "000000";
				when "010111010010" => data <= "111111";
				when "010111010011" => data <= "010010";
				when "010111010100" => data <= "010010";
				when "010111010101" => data <= "111111";
				when "010111010110" => data <= "000000";
				when "010111010111" => data <= "000000";
				when "010111011000" => data <= "000000";
				when "010111011001" => data <= "000000";
				when "010111011010" => data <= "000000";
				when "010111011011" => data <= "111111";
				when "010111011100" => data <= "010010";
				when "010111011101" => data <= "010010";
				when "010111011110" => data <= "111111";
				when "010111011111" => data <= "000000";
				when "010111100000" => data <= "000000";
				when "010111100001" => data <= "000000";
				when "010111100010" => data <= "000000";
				when "010111100011" => data <= "000000";
				when "010111100100" => data <= "000000";
				when "010111100101" => data <= "111111";
				when "010111100110" => data <= "010010";
				when "010111100111" => data <= "010010";
				when "010111101000" => data <= "111111";
				when "010111101001" => data <= "000000";
				when "010111101010" => data <= "000000";
				when "010111101011" => data <= "000000";
				when "010111101100" => data <= "000000";
				when "010111101101" => data <= "000000";
				when "010111101110" => data <= "000000";
				when "010111101111" => data <= "000000";
				when "010111110000" => data <= "000000";
				when "010111110001" => data <= "000000";
				when "010111110010" => data <= "000000";
				when "010111110011" => data <= "000000";
				when "010111110100" => data <= "000000";
				when "010111110101" => data <= "000000";
				when "010111110110" => data <= "000000";
				when "010111110111" => data <= "000000";
				when "010111111000" => data <= "000000";
				when "010111111001" => data <= "000000";
				when "010111111010" => data <= "000000";
				when "010111111011" => data <= "000000";
				when "010111111100" => data <= "000000";
				when "010111111101" => data <= "000000";
				when "010111111110" => data <= "000000";
				when "010111111111" => data <= "000000";
				when "011000000000" => data <= "000000";
				when "011000000001" => data <= "000000";
				when "011000000010" => data <= "000000";
				when "011000000011" => data <= "000000";
				when "011000000100" => data <= "000000";
				when "011000000101" => data <= "000000";
				when "011000000110" => data <= "000000";
				when "011000000111" => data <= "000000";
				when "011000001000" => data <= "000000";
				when "011000001001" => data <= "000000";
				when "011000001010" => data <= "000000";
				when "011000001011" => data <= "000000";
				when "011000001100" => data <= "000000";
				when "011000001101" => data <= "000000";
				when "011000001110" => data <= "000000";
				when "011000001111" => data <= "000000";
				when "011000010000" => data <= "000000";
				when "011000010001" => data <= "000000";
				when "011000010010" => data <= "000000";
				when "011000010011" => data <= "000000";
				when "011000010100" => data <= "111111";
				when "011000010101" => data <= "010011";
				when "011000010110" => data <= "010011";
				when "011000010111" => data <= "111111";
				when "011000011000" => data <= "000000";
				when "011000011001" => data <= "000000";
				when "011000011010" => data <= "000000";
				when "011000011011" => data <= "000000";
				when "011000011100" => data <= "111111";
				when "011000011101" => data <= "010011";
				when "011000011110" => data <= "010011";
				when "011000011111" => data <= "111111";
				when "011000100000" => data <= "000000";
				when "011000100001" => data <= "000000";
				when "011000100010" => data <= "000000";
				when "011000100011" => data <= "000000";
				when "011000100100" => data <= "000000";
				when "011000100101" => data <= "000000";
				when "011000100110" => data <= "111111";
				when "011000100111" => data <= "010011";
				when "011000101000" => data <= "010011";
				when "011000101001" => data <= "111111";
				when "011000101010" => data <= "000000";
				when "011000101011" => data <= "000000";
				when "011000101100" => data <= "000000";
				when "011000101101" => data <= "000000";
				when "011000101110" => data <= "000000";
				when "011000101111" => data <= "000000";
				when "011000110000" => data <= "000000";
				when "011000110001" => data <= "000000";
				when "011000110010" => data <= "000000";
				when "011000110011" => data <= "000000";
				when "011000110100" => data <= "000000";
				when "011000110101" => data <= "000000";
				when "011000110110" => data <= "000000";
				when "011000110111" => data <= "000000";
				when "011000111000" => data <= "000000";
				when "011000111001" => data <= "000000";
				when "011000111010" => data <= "000000";
				when "011000111011" => data <= "000000";
				when "011000111100" => data <= "111111";
				when "011000111101" => data <= "010011";
				when "011000111110" => data <= "010011";
				when "011000111111" => data <= "111111";
				when "011001000000" => data <= "000000";
				when "011001000001" => data <= "000000";
				when "011001000010" => data <= "000000";
				when "011001000011" => data <= "000000";
				when "011001000100" => data <= "000000";
				when "011001000101" => data <= "000000";
				when "011001000110" => data <= "000000";
				when "011001000111" => data <= "000000";
				when "011001001000" => data <= "000000";
				when "011001001001" => data <= "000000";
				when "011001001010" => data <= "111111";
				when "011001001011" => data <= "010011";
				when "011001001100" => data <= "010011";
				when "011001001101" => data <= "111111";
				when "011001001110" => data <= "000000";
				when "011001001111" => data <= "000000";
				when "011001010000" => data <= "000000";
				when "011001010001" => data <= "000000";
				when "011001010010" => data <= "111111";
				when "011001010011" => data <= "010011";
				when "011001010100" => data <= "010011";
				when "011001010101" => data <= "111111";
				when "011001010110" => data <= "000000";
				when "011001010111" => data <= "000000";
				when "011001011000" => data <= "000000";
				when "011001011001" => data <= "000000";
				when "011001011010" => data <= "000000";
				when "011001011011" => data <= "111111";
				when "011001011100" => data <= "010011";
				when "011001011101" => data <= "010011";
				when "011001011110" => data <= "111111";
				when "011001011111" => data <= "000000";
				when "011001100000" => data <= "000000";
				when "011001100001" => data <= "000000";
				when "011001100010" => data <= "000000";
				when "011001100011" => data <= "000000";
				when "011001100100" => data <= "000000";
				when "011001100101" => data <= "111111";
				when "011001100110" => data <= "010011";
				when "011001100111" => data <= "010011";
				when "011001101000" => data <= "111111";
				when "011001101001" => data <= "000000";
				when "011001101010" => data <= "000000";
				when "011001101011" => data <= "000000";
				when "011001101100" => data <= "000000";
				when "011001101101" => data <= "000000";
				when "011001101110" => data <= "000000";
				when "011001101111" => data <= "000000";
				when "011001110000" => data <= "000000";
				when "011001110001" => data <= "000000";
				when "011001110010" => data <= "000000";
				when "011001110011" => data <= "000000";
				when "011001110100" => data <= "000000";
				when "011001110101" => data <= "000000";
				when "011001110110" => data <= "000000";
				when "011001110111" => data <= "000000";
				when "011001111000" => data <= "000000";
				when "011001111001" => data <= "000000";
				when "011001111010" => data <= "000000";
				when "011001111011" => data <= "000000";
				when "011001111100" => data <= "000000";
				when "011001111101" => data <= "000000";
				when "011001111110" => data <= "000000";
				when "011001111111" => data <= "000000";
				when "011010000000" => data <= "000000";
				when "011010000001" => data <= "000000";
				when "011010000010" => data <= "000000";
				when "011010000011" => data <= "000000";
				when "011010000100" => data <= "000000";
				when "011010000101" => data <= "000000";
				when "011010000110" => data <= "000000";
				when "011010000111" => data <= "000000";
				when "011010001000" => data <= "000000";
				when "011010001001" => data <= "000000";
				when "011010001010" => data <= "000000";
				when "011010001011" => data <= "000000";
				when "011010001100" => data <= "000000";
				when "011010001101" => data <= "000000";
				when "011010001110" => data <= "000000";
				when "011010001111" => data <= "000000";
				when "011010010000" => data <= "000000";
				when "011010010001" => data <= "000000";
				when "011010010010" => data <= "000000";
				when "011010010011" => data <= "000000";
				when "011010010100" => data <= "111111";
				when "011010010101" => data <= "010011";
				when "011010010110" => data <= "010011";
				when "011010010111" => data <= "111111";
				when "011010011000" => data <= "000000";
				when "011010011001" => data <= "000000";
				when "011010011010" => data <= "000000";
				when "011010011011" => data <= "000000";
				when "011010011100" => data <= "111111";
				when "011010011101" => data <= "010011";
				when "011010011110" => data <= "010011";
				when "011010011111" => data <= "111111";
				when "011010100000" => data <= "000000";
				when "011010100001" => data <= "000000";
				when "011010100010" => data <= "000000";
				when "011010100011" => data <= "000000";
				when "011010100100" => data <= "000000";
				when "011010100101" => data <= "000000";
				when "011010100110" => data <= "111111";
				when "011010100111" => data <= "010011";
				when "011010101000" => data <= "010011";
				when "011010101001" => data <= "111111";
				when "011010101010" => data <= "000000";
				when "011010101011" => data <= "000000";
				when "011010101100" => data <= "000000";
				when "011010101101" => data <= "000000";
				when "011010101110" => data <= "000000";
				when "011010101111" => data <= "000000";
				when "011010110000" => data <= "000000";
				when "011010110001" => data <= "000000";
				when "011010110010" => data <= "000000";
				when "011010110011" => data <= "000000";
				when "011010110100" => data <= "000000";
				when "011010110101" => data <= "000000";
				when "011010110110" => data <= "000000";
				when "011010110111" => data <= "000000";
				when "011010111000" => data <= "000000";
				when "011010111001" => data <= "000000";
				when "011010111010" => data <= "000000";
				when "011010111011" => data <= "000000";
				when "011010111100" => data <= "111111";
				when "011010111101" => data <= "010011";
				when "011010111110" => data <= "010011";
				when "011010111111" => data <= "111111";
				when "011011000000" => data <= "000000";
				when "011011000001" => data <= "000000";
				when "011011000010" => data <= "000000";
				when "011011000011" => data <= "000000";
				when "011011000100" => data <= "000000";
				when "011011000101" => data <= "000000";
				when "011011000110" => data <= "000000";
				when "011011000111" => data <= "000000";
				when "011011001000" => data <= "000000";
				when "011011001001" => data <= "000000";
				when "011011001010" => data <= "111111";
				when "011011001011" => data <= "010011";
				when "011011001100" => data <= "010011";
				when "011011001101" => data <= "111111";
				when "011011001110" => data <= "000000";
				when "011011001111" => data <= "000000";
				when "011011010000" => data <= "000000";
				when "011011010001" => data <= "000000";
				when "011011010010" => data <= "111111";
				when "011011010011" => data <= "010011";
				when "011011010100" => data <= "010011";
				when "011011010101" => data <= "111111";
				when "011011010110" => data <= "000000";
				when "011011010111" => data <= "000000";
				when "011011011000" => data <= "000000";
				when "011011011001" => data <= "000000";
				when "011011011010" => data <= "000000";
				when "011011011011" => data <= "111111";
				when "011011011100" => data <= "010011";
				when "011011011101" => data <= "010011";
				when "011011011110" => data <= "111111";
				when "011011011111" => data <= "000000";
				when "011011100000" => data <= "000000";
				when "011011100001" => data <= "000000";
				when "011011100010" => data <= "000000";
				when "011011100011" => data <= "000000";
				when "011011100100" => data <= "000000";
				when "011011100101" => data <= "111111";
				when "011011100110" => data <= "010011";
				when "011011100111" => data <= "010011";
				when "011011101000" => data <= "111111";
				when "011011101001" => data <= "000000";
				when "011011101010" => data <= "000000";
				when "011011101011" => data <= "000000";
				when "011011101100" => data <= "000000";
				when "011011101101" => data <= "000000";
				when "011011101110" => data <= "000000";
				when "011011101111" => data <= "000000";
				when "011011110000" => data <= "000000";
				when "011011110001" => data <= "000000";
				when "011011110010" => data <= "000000";
				when "011011110011" => data <= "000000";
				when "011011110100" => data <= "000000";
				when "011011110101" => data <= "000000";
				when "011011110110" => data <= "000000";
				when "011011110111" => data <= "000000";
				when "011011111000" => data <= "000000";
				when "011011111001" => data <= "000000";
				when "011011111010" => data <= "000000";
				when "011011111011" => data <= "000000";
				when "011011111100" => data <= "000000";
				when "011011111101" => data <= "000000";
				when "011011111110" => data <= "000000";
				when "011011111111" => data <= "000000";
				when "011100000000" => data <= "000000";
				when "011100000001" => data <= "000000";
				when "011100000010" => data <= "000000";
				when "011100000011" => data <= "000000";
				when "011100000100" => data <= "000000";
				when "011100000101" => data <= "000000";
				when "011100000110" => data <= "000000";
				when "011100000111" => data <= "000000";
				when "011100001000" => data <= "000000";
				when "011100001001" => data <= "000000";
				when "011100001010" => data <= "000000";
				when "011100001011" => data <= "000000";
				when "011100001100" => data <= "000000";
				when "011100001101" => data <= "000000";
				when "011100001110" => data <= "000000";
				when "011100001111" => data <= "000000";
				when "011100010000" => data <= "000000";
				when "011100010001" => data <= "000000";
				when "011100010010" => data <= "000000";
				when "011100010011" => data <= "000000";
				when "011100010100" => data <= "111111";
				when "011100010101" => data <= "010011";
				when "011100010110" => data <= "010011";
				when "011100010111" => data <= "111111";
				when "011100011000" => data <= "111111";
				when "011100011001" => data <= "111111";
				when "011100011010" => data <= "111111";
				when "011100011011" => data <= "111111";
				when "011100011100" => data <= "111111";
				when "011100011101" => data <= "010011";
				when "011100011110" => data <= "010011";
				when "011100011111" => data <= "111111";
				when "011100100000" => data <= "000000";
				when "011100100001" => data <= "000000";
				when "011100100010" => data <= "000000";
				when "011100100011" => data <= "000000";
				when "011100100100" => data <= "000000";
				when "011100100101" => data <= "000000";
				when "011100100110" => data <= "111111";
				when "011100100111" => data <= "010011";
				when "011100101000" => data <= "010011";
				when "011100101001" => data <= "111111";
				when "011100101010" => data <= "111111";
				when "011100101011" => data <= "111111";
				when "011100101100" => data <= "111111";
				when "011100101101" => data <= "111111";
				when "011100101110" => data <= "111111";
				when "011100101111" => data <= "000000";
				when "011100110000" => data <= "000000";
				when "011100110001" => data <= "000000";
				when "011100110010" => data <= "000000";
				when "011100110011" => data <= "000000";
				when "011100110100" => data <= "000000";
				when "011100110101" => data <= "000000";
				when "011100110110" => data <= "000000";
				when "011100110111" => data <= "000000";
				when "011100111000" => data <= "000000";
				when "011100111001" => data <= "000000";
				when "011100111010" => data <= "000000";
				when "011100111011" => data <= "000000";
				when "011100111100" => data <= "111111";
				when "011100111101" => data <= "010011";
				when "011100111110" => data <= "010011";
				when "011100111111" => data <= "111111";
				when "011101000000" => data <= "000000";
				when "011101000001" => data <= "000000";
				when "011101000010" => data <= "000000";
				when "011101000011" => data <= "000000";
				when "011101000100" => data <= "000000";
				when "011101000101" => data <= "000000";
				when "011101000110" => data <= "000000";
				when "011101000111" => data <= "000000";
				when "011101001000" => data <= "000000";
				when "011101001001" => data <= "000000";
				when "011101001010" => data <= "111111";
				when "011101001011" => data <= "010011";
				when "011101001100" => data <= "010011";
				when "011101001101" => data <= "111111";
				when "011101001110" => data <= "111111";
				when "011101001111" => data <= "111111";
				when "011101010000" => data <= "111111";
				when "011101010001" => data <= "111111";
				when "011101010010" => data <= "111111";
				when "011101010011" => data <= "010011";
				when "011101010100" => data <= "010011";
				when "011101010101" => data <= "111111";
				when "011101010110" => data <= "000000";
				when "011101010111" => data <= "000000";
				when "011101011000" => data <= "000000";
				when "011101011001" => data <= "000000";
				when "011101011010" => data <= "000000";
				when "011101011011" => data <= "111111";
				when "011101011100" => data <= "010011";
				when "011101011101" => data <= "010011";
				when "011101011110" => data <= "111111";
				when "011101011111" => data <= "000000";
				when "011101100000" => data <= "000000";
				when "011101100001" => data <= "000000";
				when "011101100010" => data <= "000000";
				when "011101100011" => data <= "000000";
				when "011101100100" => data <= "000000";
				when "011101100101" => data <= "111111";
				when "011101100110" => data <= "010011";
				when "011101100111" => data <= "010011";
				when "011101101000" => data <= "111111";
				when "011101101001" => data <= "000000";
				when "011101101010" => data <= "000000";
				when "011101101011" => data <= "000000";
				when "011101101100" => data <= "000000";
				when "011101101101" => data <= "000000";
				when "011101101110" => data <= "000000";
				when "011101101111" => data <= "000000";
				when "011101110000" => data <= "000000";
				when "011101110001" => data <= "000000";
				when "011101110010" => data <= "000000";
				when "011101110011" => data <= "000000";
				when "011101110100" => data <= "000000";
				when "011101110101" => data <= "000000";
				when "011101110110" => data <= "000000";
				when "011101110111" => data <= "000000";
				when "011101111000" => data <= "000000";
				when "011101111001" => data <= "000000";
				when "011101111010" => data <= "000000";
				when "011101111011" => data <= "000000";
				when "011101111100" => data <= "000000";
				when "011101111101" => data <= "000000";
				when "011101111110" => data <= "000000";
				when "011101111111" => data <= "000000";
				when "011110000000" => data <= "000000";
				when "011110000001" => data <= "000000";
				when "011110000010" => data <= "000000";
				when "011110000011" => data <= "000000";
				when "011110000100" => data <= "000000";
				when "011110000101" => data <= "000000";
				when "011110000110" => data <= "000000";
				when "011110000111" => data <= "000000";
				when "011110001000" => data <= "000000";
				when "011110001001" => data <= "000000";
				when "011110001010" => data <= "000000";
				when "011110001011" => data <= "000000";
				when "011110001100" => data <= "000000";
				when "011110001101" => data <= "000000";
				when "011110001110" => data <= "000000";
				when "011110001111" => data <= "000000";
				when "011110010000" => data <= "000000";
				when "011110010001" => data <= "000000";
				when "011110010010" => data <= "000000";
				when "011110010011" => data <= "000000";
				when "011110010100" => data <= "111111";
				when "011110010101" => data <= "010011";
				when "011110010110" => data <= "010011";
				when "011110010111" => data <= "010011";
				when "011110011000" => data <= "010011";
				when "011110011001" => data <= "010011";
				when "011110011010" => data <= "010011";
				when "011110011011" => data <= "010011";
				when "011110011100" => data <= "010011";
				when "011110011101" => data <= "111111";
				when "011110011110" => data <= "111111";
				when "011110011111" => data <= "000000";
				when "011110100000" => data <= "000000";
				when "011110100001" => data <= "000000";
				when "011110100010" => data <= "000000";
				when "011110100011" => data <= "000000";
				when "011110100100" => data <= "000000";
				when "011110100101" => data <= "000000";
				when "011110100110" => data <= "111111";
				when "011110100111" => data <= "010011";
				when "011110101000" => data <= "010011";
				when "011110101001" => data <= "010011";
				when "011110101010" => data <= "010011";
				when "011110101011" => data <= "010011";
				when "011110101100" => data <= "010011";
				when "011110101101" => data <= "010011";
				when "011110101110" => data <= "010011";
				when "011110101111" => data <= "111111";
				when "011110110000" => data <= "000000";
				when "011110110001" => data <= "000000";
				when "011110110010" => data <= "000000";
				when "011110110011" => data <= "000000";
				when "011110110100" => data <= "000000";
				when "011110110101" => data <= "000000";
				when "011110110110" => data <= "000000";
				when "011110110111" => data <= "000000";
				when "011110111000" => data <= "000000";
				when "011110111001" => data <= "000000";
				when "011110111010" => data <= "000000";
				when "011110111011" => data <= "000000";
				when "011110111100" => data <= "111111";
				when "011110111101" => data <= "010011";
				when "011110111110" => data <= "010011";
				when "011110111111" => data <= "111111";
				when "011111000000" => data <= "000000";
				when "011111000001" => data <= "000000";
				when "011111000010" => data <= "000000";
				when "011111000011" => data <= "000000";
				when "011111000100" => data <= "000000";
				when "011111000101" => data <= "000000";
				when "011111000110" => data <= "000000";
				when "011111000111" => data <= "000000";
				when "011111001000" => data <= "000000";
				when "011111001001" => data <= "000000";
				when "011111001010" => data <= "111111";
				when "011111001011" => data <= "010011";
				when "011111001100" => data <= "010011";
				when "011111001101" => data <= "010011";
				when "011111001110" => data <= "010011";
				when "011111001111" => data <= "010011";
				when "011111010000" => data <= "010011";
				when "011111010001" => data <= "010011";
				when "011111010010" => data <= "010011";
				when "011111010011" => data <= "111111";
				when "011111010100" => data <= "111111";
				when "011111010101" => data <= "000000";
				when "011111010110" => data <= "000000";
				when "011111010111" => data <= "000000";
				when "011111011000" => data <= "000000";
				when "011111011001" => data <= "000000";
				when "011111011010" => data <= "000000";
				when "011111011011" => data <= "111111";
				when "011111011100" => data <= "010011";
				when "011111011101" => data <= "010011";
				when "011111011110" => data <= "111111";
				when "011111011111" => data <= "000000";
				when "011111100000" => data <= "000000";
				when "011111100001" => data <= "000000";
				when "011111100010" => data <= "000000";
				when "011111100011" => data <= "000000";
				when "011111100100" => data <= "000000";
				when "011111100101" => data <= "111111";
				when "011111100110" => data <= "010011";
				when "011111100111" => data <= "010011";
				when "011111101000" => data <= "111111";
				when "011111101001" => data <= "000000";
				when "011111101010" => data <= "000000";
				when "011111101011" => data <= "000000";
				when "011111101100" => data <= "000000";
				when "011111101101" => data <= "000000";
				when "011111101110" => data <= "000000";
				when "011111101111" => data <= "000000";
				when "011111110000" => data <= "000000";
				when "011111110001" => data <= "000000";
				when "011111110010" => data <= "000000";
				when "011111110011" => data <= "000000";
				when "011111110100" => data <= "000000";
				when "011111110101" => data <= "000000";
				when "011111110110" => data <= "000000";
				when "011111110111" => data <= "000000";
				when "011111111000" => data <= "000000";
				when "011111111001" => data <= "000000";
				when "011111111010" => data <= "000000";
				when "011111111011" => data <= "000000";
				when "011111111100" => data <= "000000";
				when "011111111101" => data <= "000000";
				when "011111111110" => data <= "000000";
				when "011111111111" => data <= "000000";
				when "100000000000" => data <= "000000";
				when "100000000001" => data <= "000000";
				when "100000000010" => data <= "000000";
				when "100000000011" => data <= "000000";
				when "100000000100" => data <= "000000";
				when "100000000101" => data <= "000000";
				when "100000000110" => data <= "000000";
				when "100000000111" => data <= "000000";
				when "100000001000" => data <= "000000";
				when "100000001001" => data <= "000000";
				when "100000001010" => data <= "000000";
				when "100000001011" => data <= "000000";
				when "100000001100" => data <= "000000";
				when "100000001101" => data <= "000000";
				when "100000001110" => data <= "000000";
				when "100000001111" => data <= "000000";
				when "100000010000" => data <= "000000";
				when "100000010001" => data <= "000000";
				when "100000010010" => data <= "000000";
				when "100000010011" => data <= "000000";
				when "100000010100" => data <= "111111";
				when "100000010101" => data <= "010011";
				when "100000010110" => data <= "010011";
				when "100000010111" => data <= "010011";
				when "100000011000" => data <= "010011";
				when "100000011001" => data <= "010011";
				when "100000011010" => data <= "010011";
				when "100000011011" => data <= "010011";
				when "100000011100" => data <= "010011";
				when "100000011101" => data <= "111111";
				when "100000011110" => data <= "000000";
				when "100000011111" => data <= "000000";
				when "100000100000" => data <= "000000";
				when "100000100001" => data <= "000000";
				when "100000100010" => data <= "000000";
				when "100000100011" => data <= "000000";
				when "100000100100" => data <= "000000";
				when "100000100101" => data <= "000000";
				when "100000100110" => data <= "111111";
				when "100000100111" => data <= "010011";
				when "100000101000" => data <= "010011";
				when "100000101001" => data <= "010011";
				when "100000101010" => data <= "010011";
				when "100000101011" => data <= "010011";
				when "100000101100" => data <= "010011";
				when "100000101101" => data <= "010011";
				when "100000101110" => data <= "010011";
				when "100000101111" => data <= "111111";
				when "100000110000" => data <= "000000";
				when "100000110001" => data <= "000000";
				when "100000110010" => data <= "000000";
				when "100000110011" => data <= "000000";
				when "100000110100" => data <= "000000";
				when "100000110101" => data <= "000000";
				when "100000110110" => data <= "000000";
				when "100000110111" => data <= "000000";
				when "100000111000" => data <= "000000";
				when "100000111001" => data <= "000000";
				when "100000111010" => data <= "000000";
				when "100000111011" => data <= "000000";
				when "100000111100" => data <= "111111";
				when "100000111101" => data <= "100011";
				when "100000111110" => data <= "100011";
				when "100000111111" => data <= "111111";
				when "100001000000" => data <= "000000";
				when "100001000001" => data <= "000000";
				when "100001000010" => data <= "000000";
				when "100001000011" => data <= "000000";
				when "100001000100" => data <= "000000";
				when "100001000101" => data <= "000000";
				when "100001000110" => data <= "000000";
				when "100001000111" => data <= "000000";
				when "100001001000" => data <= "000000";
				when "100001001001" => data <= "000000";
				when "100001001010" => data <= "111111";
				when "100001001011" => data <= "100011";
				when "100001001100" => data <= "100011";
				when "100001001101" => data <= "010011";
				when "100001001110" => data <= "010011";
				when "100001001111" => data <= "010011";
				when "100001010000" => data <= "010011";
				when "100001010001" => data <= "010011";
				when "100001010010" => data <= "010011";
				when "100001010011" => data <= "111111";
				when "100001010100" => data <= "000000";
				when "100001010101" => data <= "000000";
				when "100001010110" => data <= "000000";
				when "100001010111" => data <= "000000";
				when "100001011000" => data <= "000000";
				when "100001011001" => data <= "000000";
				when "100001011010" => data <= "000000";
				when "100001011011" => data <= "111111";
				when "100001011100" => data <= "100011";
				when "100001011101" => data <= "100011";
				when "100001011110" => data <= "111111";
				when "100001011111" => data <= "000000";
				when "100001100000" => data <= "000000";
				when "100001100001" => data <= "000000";
				when "100001100010" => data <= "000000";
				when "100001100011" => data <= "000000";
				when "100001100100" => data <= "000000";
				when "100001100101" => data <= "111111";
				when "100001100110" => data <= "100011";
				when "100001100111" => data <= "100011";
				when "100001101000" => data <= "111111";
				when "100001101001" => data <= "000000";
				when "100001101010" => data <= "000000";
				when "100001101011" => data <= "000000";
				when "100001101100" => data <= "000000";
				when "100001101101" => data <= "000000";
				when "100001101110" => data <= "000000";
				when "100001101111" => data <= "000000";
				when "100001110000" => data <= "000000";
				when "100001110001" => data <= "000000";
				when "100001110010" => data <= "000000";
				when "100001110011" => data <= "000000";
				when "100001110100" => data <= "000000";
				when "100001110101" => data <= "000000";
				when "100001110110" => data <= "000000";
				when "100001110111" => data <= "000000";
				when "100001111000" => data <= "000000";
				when "100001111001" => data <= "000000";
				when "100001111010" => data <= "000000";
				when "100001111011" => data <= "000000";
				when "100001111100" => data <= "000000";
				when "100001111101" => data <= "000000";
				when "100001111110" => data <= "000000";
				when "100001111111" => data <= "000000";
				when "100010000000" => data <= "000000";
				when "100010000001" => data <= "000000";
				when "100010000010" => data <= "000000";
				when "100010000011" => data <= "000000";
				when "100010000100" => data <= "000000";
				when "100010000101" => data <= "000000";
				when "100010000110" => data <= "000000";
				when "100010000111" => data <= "000000";
				when "100010001000" => data <= "000000";
				when "100010001001" => data <= "000000";
				when "100010001010" => data <= "000000";
				when "100010001011" => data <= "000000";
				when "100010001100" => data <= "000000";
				when "100010001101" => data <= "000000";
				when "100010001110" => data <= "000000";
				when "100010001111" => data <= "000000";
				when "100010010000" => data <= "000000";
				when "100010010001" => data <= "000000";
				when "100010010010" => data <= "000000";
				when "100010010011" => data <= "000000";
				when "100010010100" => data <= "111111";
				when "100010010101" => data <= "100011";
				when "100010010110" => data <= "100011";
				when "100010010111" => data <= "111111";
				when "100010011000" => data <= "111111";
				when "100010011001" => data <= "111111";
				when "100010011010" => data <= "111111";
				when "100010011011" => data <= "111111";
				when "100010011100" => data <= "111111";
				when "100010011101" => data <= "100011";
				when "100010011110" => data <= "111111";
				when "100010011111" => data <= "000000";
				when "100010100000" => data <= "000000";
				when "100010100001" => data <= "000000";
				when "100010100010" => data <= "000000";
				when "100010100011" => data <= "000000";
				when "100010100100" => data <= "000000";
				when "100010100101" => data <= "000000";
				when "100010100110" => data <= "111111";
				when "100010100111" => data <= "100011";
				when "100010101000" => data <= "100011";
				when "100010101001" => data <= "111111";
				when "100010101010" => data <= "111111";
				when "100010101011" => data <= "111111";
				when "100010101100" => data <= "111111";
				when "100010101101" => data <= "111111";
				when "100010101110" => data <= "111111";
				when "100010101111" => data <= "000000";
				when "100010110000" => data <= "000000";
				when "100010110001" => data <= "000000";
				when "100010110010" => data <= "000000";
				when "100010110011" => data <= "000000";
				when "100010110100" => data <= "000000";
				when "100010110101" => data <= "000000";
				when "100010110110" => data <= "000000";
				when "100010110111" => data <= "000000";
				when "100010111000" => data <= "000000";
				when "100010111001" => data <= "000000";
				when "100010111010" => data <= "000000";
				when "100010111011" => data <= "000000";
				when "100010111100" => data <= "111111";
				when "100010111101" => data <= "100011";
				when "100010111110" => data <= "100011";
				when "100010111111" => data <= "111111";
				when "100011000000" => data <= "000000";
				when "100011000001" => data <= "000000";
				when "100011000010" => data <= "000000";
				when "100011000011" => data <= "000000";
				when "100011000100" => data <= "000000";
				when "100011000101" => data <= "000000";
				when "100011000110" => data <= "000000";
				when "100011000111" => data <= "000000";
				when "100011001000" => data <= "000000";
				when "100011001001" => data <= "000000";
				when "100011001010" => data <= "111111";
				when "100011001011" => data <= "100011";
				when "100011001100" => data <= "100011";
				when "100011001101" => data <= "111111";
				when "100011001110" => data <= "111111";
				when "100011001111" => data <= "111111";
				when "100011010000" => data <= "111111";
				when "100011010001" => data <= "111111";
				when "100011010010" => data <= "111111";
				when "100011010011" => data <= "100011";
				when "100011010100" => data <= "111111";
				when "100011010101" => data <= "000000";
				when "100011010110" => data <= "000000";
				when "100011010111" => data <= "000000";
				when "100011011000" => data <= "000000";
				when "100011011001" => data <= "000000";
				when "100011011010" => data <= "000000";
				when "100011011011" => data <= "111111";
				when "100011011100" => data <= "100011";
				when "100011011101" => data <= "100011";
				when "100011011110" => data <= "111111";
				when "100011011111" => data <= "000000";
				when "100011100000" => data <= "000000";
				when "100011100001" => data <= "000000";
				when "100011100010" => data <= "000000";
				when "100011100011" => data <= "000000";
				when "100011100100" => data <= "000000";
				when "100011100101" => data <= "111111";
				when "100011100110" => data <= "100011";
				when "100011100111" => data <= "100011";
				when "100011101000" => data <= "111111";
				when "100011101001" => data <= "000000";
				when "100011101010" => data <= "000000";
				when "100011101011" => data <= "000000";
				when "100011101100" => data <= "000000";
				when "100011101101" => data <= "000000";
				when "100011101110" => data <= "000000";
				when "100011101111" => data <= "000000";
				when "100011110000" => data <= "000000";
				when "100011110001" => data <= "000000";
				when "100011110010" => data <= "000000";
				when "100011110011" => data <= "000000";
				when "100011110100" => data <= "000000";
				when "100011110101" => data <= "000000";
				when "100011110110" => data <= "000000";
				when "100011110111" => data <= "000000";
				when "100011111000" => data <= "000000";
				when "100011111001" => data <= "000000";
				when "100011111010" => data <= "000000";
				when "100011111011" => data <= "000000";
				when "100011111100" => data <= "000000";
				when "100011111101" => data <= "000000";
				when "100011111110" => data <= "000000";
				when "100011111111" => data <= "000000";
				when "100100000000" => data <= "000000";
				when "100100000001" => data <= "000000";
				when "100100000010" => data <= "000000";
				when "100100000011" => data <= "000000";
				when "100100000100" => data <= "000000";
				when "100100000101" => data <= "000000";
				when "100100000110" => data <= "000000";
				when "100100000111" => data <= "000000";
				when "100100001000" => data <= "000000";
				when "100100001001" => data <= "000000";
				when "100100001010" => data <= "000000";
				when "100100001011" => data <= "000000";
				when "100100001100" => data <= "000000";
				when "100100001101" => data <= "000000";
				when "100100001110" => data <= "000000";
				when "100100001111" => data <= "000000";
				when "100100010000" => data <= "000000";
				when "100100010001" => data <= "000000";
				when "100100010010" => data <= "000000";
				when "100100010011" => data <= "000000";
				when "100100010100" => data <= "111111";
				when "100100010101" => data <= "100011";
				when "100100010110" => data <= "100011";
				when "100100010111" => data <= "111111";
				when "100100011000" => data <= "000000";
				when "100100011001" => data <= "000000";
				when "100100011010" => data <= "000000";
				when "100100011011" => data <= "000000";
				when "100100011100" => data <= "111111";
				when "100100011101" => data <= "100011";
				when "100100011110" => data <= "100011";
				when "100100011111" => data <= "111111";
				when "100100100000" => data <= "000000";
				when "100100100001" => data <= "000000";
				when "100100100010" => data <= "000000";
				when "100100100011" => data <= "000000";
				when "100100100100" => data <= "000000";
				when "100100100101" => data <= "000000";
				when "100100100110" => data <= "111111";
				when "100100100111" => data <= "100011";
				when "100100101000" => data <= "100011";
				when "100100101001" => data <= "111111";
				when "100100101010" => data <= "000000";
				when "100100101011" => data <= "000000";
				when "100100101100" => data <= "000000";
				when "100100101101" => data <= "000000";
				when "100100101110" => data <= "000000";
				when "100100101111" => data <= "000000";
				when "100100110000" => data <= "000000";
				when "100100110001" => data <= "000000";
				when "100100110010" => data <= "000000";
				when "100100110011" => data <= "000000";
				when "100100110100" => data <= "000000";
				when "100100110101" => data <= "000000";
				when "100100110110" => data <= "000000";
				when "100100110111" => data <= "000000";
				when "100100111000" => data <= "000000";
				when "100100111001" => data <= "000000";
				when "100100111010" => data <= "000000";
				when "100100111011" => data <= "000000";
				when "100100111100" => data <= "111111";
				when "100100111101" => data <= "100011";
				when "100100111110" => data <= "100011";
				when "100100111111" => data <= "111111";
				when "100101000000" => data <= "000000";
				when "100101000001" => data <= "000000";
				when "100101000010" => data <= "000000";
				when "100101000011" => data <= "000000";
				when "100101000100" => data <= "000000";
				when "100101000101" => data <= "000000";
				when "100101000110" => data <= "000000";
				when "100101000111" => data <= "000000";
				when "100101001000" => data <= "000000";
				when "100101001001" => data <= "000000";
				when "100101001010" => data <= "111111";
				when "100101001011" => data <= "100011";
				when "100101001100" => data <= "100011";
				when "100101001101" => data <= "111111";
				when "100101001110" => data <= "000000";
				when "100101001111" => data <= "000000";
				when "100101010000" => data <= "000000";
				when "100101010001" => data <= "000000";
				when "100101010010" => data <= "111111";
				when "100101010011" => data <= "100011";
				when "100101010100" => data <= "100011";
				when "100101010101" => data <= "111111";
				when "100101010110" => data <= "000000";
				when "100101010111" => data <= "000000";
				when "100101011000" => data <= "000000";
				when "100101011001" => data <= "000000";
				when "100101011010" => data <= "000000";
				when "100101011011" => data <= "111111";
				when "100101011100" => data <= "100011";
				when "100101011101" => data <= "100011";
				when "100101011110" => data <= "111111";
				when "100101011111" => data <= "000000";
				when "100101100000" => data <= "000000";
				when "100101100001" => data <= "000000";
				when "100101100010" => data <= "000000";
				when "100101100011" => data <= "000000";
				when "100101100100" => data <= "000000";
				when "100101100101" => data <= "111111";
				when "100101100110" => data <= "100011";
				when "100101100111" => data <= "100011";
				when "100101101000" => data <= "111111";
				when "100101101001" => data <= "000000";
				when "100101101010" => data <= "000000";
				when "100101101011" => data <= "000000";
				when "100101101100" => data <= "000000";
				when "100101101101" => data <= "000000";
				when "100101101110" => data <= "000000";
				when "100101101111" => data <= "000000";
				when "100101110000" => data <= "000000";
				when "100101110001" => data <= "000000";
				when "100101110010" => data <= "000000";
				when "100101110011" => data <= "000000";
				when "100101110100" => data <= "000000";
				when "100101110101" => data <= "000000";
				when "100101110110" => data <= "000000";
				when "100101110111" => data <= "000000";
				when "100101111000" => data <= "000000";
				when "100101111001" => data <= "000000";
				when "100101111010" => data <= "000000";
				when "100101111011" => data <= "000000";
				when "100101111100" => data <= "000000";
				when "100101111101" => data <= "000000";
				when "100101111110" => data <= "000000";
				when "100101111111" => data <= "000000";
				when "100110000000" => data <= "000000";
				when "100110000001" => data <= "000000";
				when "100110000010" => data <= "000000";
				when "100110000011" => data <= "000000";
				when "100110000100" => data <= "000000";
				when "100110000101" => data <= "000000";
				when "100110000110" => data <= "000000";
				when "100110000111" => data <= "000000";
				when "100110001000" => data <= "000000";
				when "100110001001" => data <= "000000";
				when "100110001010" => data <= "000000";
				when "100110001011" => data <= "000000";
				when "100110001100" => data <= "000000";
				when "100110001101" => data <= "000000";
				when "100110001110" => data <= "000000";
				when "100110001111" => data <= "000000";
				when "100110010000" => data <= "000000";
				when "100110010001" => data <= "000000";
				when "100110010010" => data <= "000000";
				when "100110010011" => data <= "000000";
				when "100110010100" => data <= "111111";
				when "100110010101" => data <= "100011";
				when "100110010110" => data <= "100011";
				when "100110010111" => data <= "111111";
				when "100110011000" => data <= "000000";
				when "100110011001" => data <= "000000";
				when "100110011010" => data <= "000000";
				when "100110011011" => data <= "000000";
				when "100110011100" => data <= "111111";
				when "100110011101" => data <= "100011";
				when "100110011110" => data <= "100011";
				when "100110011111" => data <= "111111";
				when "100110100000" => data <= "000000";
				when "100110100001" => data <= "000000";
				when "100110100010" => data <= "000000";
				when "100110100011" => data <= "000000";
				when "100110100100" => data <= "000000";
				when "100110100101" => data <= "000000";
				when "100110100110" => data <= "111111";
				when "100110100111" => data <= "100011";
				when "100110101000" => data <= "100011";
				when "100110101001" => data <= "111111";
				when "100110101010" => data <= "000000";
				when "100110101011" => data <= "000000";
				when "100110101100" => data <= "000000";
				when "100110101101" => data <= "000000";
				when "100110101110" => data <= "000000";
				when "100110101111" => data <= "000000";
				when "100110110000" => data <= "000000";
				when "100110110001" => data <= "000000";
				when "100110110010" => data <= "000000";
				when "100110110011" => data <= "000000";
				when "100110110100" => data <= "000000";
				when "100110110101" => data <= "000000";
				when "100110110110" => data <= "000000";
				when "100110110111" => data <= "000000";
				when "100110111000" => data <= "000000";
				when "100110111001" => data <= "000000";
				when "100110111010" => data <= "000000";
				when "100110111011" => data <= "000000";
				when "100110111100" => data <= "111111";
				when "100110111101" => data <= "100011";
				when "100110111110" => data <= "100011";
				when "100110111111" => data <= "111111";
				when "100111000000" => data <= "000000";
				when "100111000001" => data <= "000000";
				when "100111000010" => data <= "000000";
				when "100111000011" => data <= "000000";
				when "100111000100" => data <= "000000";
				when "100111000101" => data <= "000000";
				when "100111000110" => data <= "000000";
				when "100111000111" => data <= "000000";
				when "100111001000" => data <= "000000";
				when "100111001001" => data <= "000000";
				when "100111001010" => data <= "111111";
				when "100111001011" => data <= "100011";
				when "100111001100" => data <= "100011";
				when "100111001101" => data <= "111111";
				when "100111001110" => data <= "000000";
				when "100111001111" => data <= "000000";
				when "100111010000" => data <= "000000";
				when "100111010001" => data <= "000000";
				when "100111010010" => data <= "111111";
				when "100111010011" => data <= "100011";
				when "100111010100" => data <= "100011";
				when "100111010101" => data <= "111111";
				when "100111010110" => data <= "000000";
				when "100111010111" => data <= "000000";
				when "100111011000" => data <= "000000";
				when "100111011001" => data <= "000000";
				when "100111011010" => data <= "000000";
				when "100111011011" => data <= "111111";
				when "100111011100" => data <= "100011";
				when "100111011101" => data <= "100011";
				when "100111011110" => data <= "111111";
				when "100111011111" => data <= "000000";
				when "100111100000" => data <= "000000";
				when "100111100001" => data <= "000000";
				when "100111100010" => data <= "000000";
				when "100111100011" => data <= "000000";
				when "100111100100" => data <= "000000";
				when "100111100101" => data <= "111111";
				when "100111100110" => data <= "100011";
				when "100111100111" => data <= "100011";
				when "100111101000" => data <= "111111";
				when "100111101001" => data <= "000000";
				when "100111101010" => data <= "000000";
				when "100111101011" => data <= "000000";
				when "100111101100" => data <= "000000";
				when "100111101101" => data <= "000000";
				when "100111101110" => data <= "000000";
				when "100111101111" => data <= "000000";
				when "100111110000" => data <= "000000";
				when "100111110001" => data <= "000000";
				when "100111110010" => data <= "000000";
				when "100111110011" => data <= "000000";
				when "100111110100" => data <= "000000";
				when "100111110101" => data <= "000000";
				when "100111110110" => data <= "000000";
				when "100111110111" => data <= "000000";
				when "100111111000" => data <= "000000";
				when "100111111001" => data <= "000000";
				when "100111111010" => data <= "000000";
				when "100111111011" => data <= "000000";
				when "100111111100" => data <= "000000";
				when "100111111101" => data <= "000000";
				when "100111111110" => data <= "000000";
				when "100111111111" => data <= "000000";
				when "101000000000" => data <= "000000";
				when "101000000001" => data <= "000000";
				when "101000000010" => data <= "000000";
				when "101000000011" => data <= "000000";
				when "101000000100" => data <= "000000";
				when "101000000101" => data <= "000000";
				when "101000000110" => data <= "000000";
				when "101000000111" => data <= "000000";
				when "101000001000" => data <= "000000";
				when "101000001001" => data <= "000000";
				when "101000001010" => data <= "000000";
				when "101000001011" => data <= "000000";
				when "101000001100" => data <= "000000";
				when "101000001101" => data <= "000000";
				when "101000001110" => data <= "000000";
				when "101000001111" => data <= "000000";
				when "101000010000" => data <= "000000";
				when "101000010001" => data <= "000000";
				when "101000010010" => data <= "000000";
				when "101000010011" => data <= "000000";
				when "101000010100" => data <= "111111";
				when "101000010101" => data <= "100011";
				when "101000010110" => data <= "100011";
				when "101000010111" => data <= "111111";
				when "101000011000" => data <= "000000";
				when "101000011001" => data <= "000000";
				when "101000011010" => data <= "000000";
				when "101000011011" => data <= "000000";
				when "101000011100" => data <= "111111";
				when "101000011101" => data <= "100011";
				when "101000011110" => data <= "100011";
				when "101000011111" => data <= "111111";
				when "101000100000" => data <= "000000";
				when "101000100001" => data <= "000000";
				when "101000100010" => data <= "000000";
				when "101000100011" => data <= "000000";
				when "101000100100" => data <= "000000";
				when "101000100101" => data <= "000000";
				when "101000100110" => data <= "111111";
				when "101000100111" => data <= "100011";
				when "101000101000" => data <= "100011";
				when "101000101001" => data <= "111111";
				when "101000101010" => data <= "000000";
				when "101000101011" => data <= "000000";
				when "101000101100" => data <= "000000";
				when "101000101101" => data <= "000000";
				when "101000101110" => data <= "000000";
				when "101000101111" => data <= "000000";
				when "101000110000" => data <= "000000";
				when "101000110001" => data <= "000000";
				when "101000110010" => data <= "000000";
				when "101000110011" => data <= "000000";
				when "101000110100" => data <= "000000";
				when "101000110101" => data <= "000000";
				when "101000110110" => data <= "000000";
				when "101000110111" => data <= "000000";
				when "101000111000" => data <= "000000";
				when "101000111001" => data <= "000000";
				when "101000111010" => data <= "000000";
				when "101000111011" => data <= "000000";
				when "101000111100" => data <= "111111";
				when "101000111101" => data <= "100111";
				when "101000111110" => data <= "100111";
				when "101000111111" => data <= "111111";
				when "101001000000" => data <= "000000";
				when "101001000001" => data <= "000000";
				when "101001000010" => data <= "000000";
				when "101001000011" => data <= "000000";
				when "101001000100" => data <= "000000";
				when "101001000101" => data <= "000000";
				when "101001000110" => data <= "000000";
				when "101001000111" => data <= "000000";
				when "101001001000" => data <= "000000";
				when "101001001001" => data <= "000000";
				when "101001001010" => data <= "111111";
				when "101001001011" => data <= "100111";
				when "101001001100" => data <= "100111";
				when "101001001101" => data <= "111111";
				when "101001001110" => data <= "000000";
				when "101001001111" => data <= "000000";
				when "101001010000" => data <= "000000";
				when "101001010001" => data <= "000000";
				when "101001010010" => data <= "111111";
				when "101001010011" => data <= "100111";
				when "101001010100" => data <= "100111";
				when "101001010101" => data <= "111111";
				when "101001010110" => data <= "000000";
				when "101001010111" => data <= "000000";
				when "101001011000" => data <= "000000";
				when "101001011001" => data <= "000000";
				when "101001011010" => data <= "000000";
				when "101001011011" => data <= "111111";
				when "101001011100" => data <= "100111";
				when "101001011101" => data <= "100111";
				when "101001011110" => data <= "111111";
				when "101001011111" => data <= "000000";
				when "101001100000" => data <= "000000";
				when "101001100001" => data <= "000000";
				when "101001100010" => data <= "000000";
				when "101001100011" => data <= "000000";
				when "101001100100" => data <= "000000";
				when "101001100101" => data <= "111111";
				when "101001100110" => data <= "100111";
				when "101001100111" => data <= "100111";
				when "101001101000" => data <= "111111";
				when "101001101001" => data <= "000000";
				when "101001101010" => data <= "000000";
				when "101001101011" => data <= "000000";
				when "101001101100" => data <= "000000";
				when "101001101101" => data <= "000000";
				when "101001101110" => data <= "000000";
				when "101001101111" => data <= "000000";
				when "101001110000" => data <= "000000";
				when "101001110001" => data <= "000000";
				when "101001110010" => data <= "000000";
				when "101001110011" => data <= "000000";
				when "101001110100" => data <= "000000";
				when "101001110101" => data <= "000000";
				when "101001110110" => data <= "000000";
				when "101001110111" => data <= "000000";
				when "101001111000" => data <= "000000";
				when "101001111001" => data <= "000000";
				when "101001111010" => data <= "000000";
				when "101001111011" => data <= "000000";
				when "101001111100" => data <= "000000";
				when "101001111101" => data <= "000000";
				when "101001111110" => data <= "000000";
				when "101001111111" => data <= "000000";
				when "101010000000" => data <= "000000";
				when "101010000001" => data <= "000000";
				when "101010000010" => data <= "000000";
				when "101010000011" => data <= "000000";
				when "101010000100" => data <= "000000";
				when "101010000101" => data <= "000000";
				when "101010000110" => data <= "000000";
				when "101010000111" => data <= "000000";
				when "101010001000" => data <= "000000";
				when "101010001001" => data <= "000000";
				when "101010001010" => data <= "000000";
				when "101010001011" => data <= "000000";
				when "101010001100" => data <= "000000";
				when "101010001101" => data <= "000000";
				when "101010001110" => data <= "000000";
				when "101010001111" => data <= "000000";
				when "101010010000" => data <= "000000";
				when "101010010001" => data <= "000000";
				when "101010010010" => data <= "000000";
				when "101010010011" => data <= "000000";
				when "101010010100" => data <= "111111";
				when "101010010101" => data <= "100111";
				when "101010010110" => data <= "100111";
				when "101010010111" => data <= "111111";
				when "101010011000" => data <= "000000";
				when "101010011001" => data <= "000000";
				when "101010011010" => data <= "000000";
				when "101010011011" => data <= "000000";
				when "101010011100" => data <= "111111";
				when "101010011101" => data <= "100111";
				when "101010011110" => data <= "100111";
				when "101010011111" => data <= "111111";
				when "101010100000" => data <= "000000";
				when "101010100001" => data <= "000000";
				when "101010100010" => data <= "000000";
				when "101010100011" => data <= "000000";
				when "101010100100" => data <= "000000";
				when "101010100101" => data <= "000000";
				when "101010100110" => data <= "111111";
				when "101010100111" => data <= "100111";
				when "101010101000" => data <= "100111";
				when "101010101001" => data <= "111111";
				when "101010101010" => data <= "111111";
				when "101010101011" => data <= "111111";
				when "101010101100" => data <= "111111";
				when "101010101101" => data <= "111111";
				when "101010101110" => data <= "111111";
				when "101010101111" => data <= "111111";
				when "101010110000" => data <= "111111";
				when "101010110001" => data <= "000000";
				when "101010110010" => data <= "000000";
				when "101010110011" => data <= "000000";
				when "101010110100" => data <= "000000";
				when "101010110101" => data <= "000000";
				when "101010110110" => data <= "000000";
				when "101010110111" => data <= "000000";
				when "101010111000" => data <= "000000";
				when "101010111001" => data <= "000000";
				when "101010111010" => data <= "000000";
				when "101010111011" => data <= "000000";
				when "101010111100" => data <= "111111";
				when "101010111101" => data <= "100111";
				when "101010111110" => data <= "100111";
				when "101010111111" => data <= "111111";
				when "101011000000" => data <= "000000";
				when "101011000001" => data <= "000000";
				when "101011000010" => data <= "000000";
				when "101011000011" => data <= "000000";
				when "101011000100" => data <= "000000";
				when "101011000101" => data <= "000000";
				when "101011000110" => data <= "000000";
				when "101011000111" => data <= "000000";
				when "101011001000" => data <= "000000";
				when "101011001001" => data <= "000000";
				when "101011001010" => data <= "111111";
				when "101011001011" => data <= "100111";
				when "101011001100" => data <= "100111";
				when "101011001101" => data <= "111111";
				when "101011001110" => data <= "000000";
				when "101011001111" => data <= "000000";
				when "101011010000" => data <= "000000";
				when "101011010001" => data <= "000000";
				when "101011010010" => data <= "111111";
				when "101011010011" => data <= "100111";
				when "101011010100" => data <= "100111";
				when "101011010101" => data <= "111111";
				when "101011010110" => data <= "000000";
				when "101011010111" => data <= "000000";
				when "101011011000" => data <= "000000";
				when "101011011001" => data <= "000000";
				when "101011011010" => data <= "000000";
				when "101011011011" => data <= "111111";
				when "101011011100" => data <= "100111";
				when "101011011101" => data <= "100111";
				when "101011011110" => data <= "111111";
				when "101011011111" => data <= "111111";
				when "101011100000" => data <= "111111";
				when "101011100001" => data <= "111111";
				when "101011100010" => data <= "111111";
				when "101011100011" => data <= "111111";
				when "101011100100" => data <= "111111";
				when "101011100101" => data <= "111111";
				when "101011100110" => data <= "100111";
				when "101011100111" => data <= "100111";
				when "101011101000" => data <= "111111";
				when "101011101001" => data <= "000000";
				when "101011101010" => data <= "000000";
				when "101011101011" => data <= "000000";
				when "101011101100" => data <= "000000";
				when "101011101101" => data <= "000000";
				when "101011101110" => data <= "000000";
				when "101011101111" => data <= "000000";
				when "101011110000" => data <= "000000";
				when "101011110001" => data <= "000000";
				when "101011110010" => data <= "000000";
				when "101011110011" => data <= "000000";
				when "101011110100" => data <= "000000";
				when "101011110101" => data <= "000000";
				when "101011110110" => data <= "000000";
				when "101011110111" => data <= "000000";
				when "101011111000" => data <= "000000";
				when "101011111001" => data <= "000000";
				when "101011111010" => data <= "000000";
				when "101011111011" => data <= "000000";
				when "101011111100" => data <= "000000";
				when "101011111101" => data <= "000000";
				when "101011111110" => data <= "000000";
				when "101011111111" => data <= "000000";
				when "101100000000" => data <= "000000";
				when "101100000001" => data <= "000000";
				when "101100000010" => data <= "000000";
				when "101100000011" => data <= "000000";
				when "101100000100" => data <= "000000";
				when "101100000101" => data <= "000000";
				when "101100000110" => data <= "000000";
				when "101100000111" => data <= "000000";
				when "101100001000" => data <= "000000";
				when "101100001001" => data <= "000000";
				when "101100001010" => data <= "000000";
				when "101100001011" => data <= "000000";
				when "101100001100" => data <= "000000";
				when "101100001101" => data <= "000000";
				when "101100001110" => data <= "000000";
				when "101100001111" => data <= "000000";
				when "101100010000" => data <= "000000";
				when "101100010001" => data <= "000000";
				when "101100010010" => data <= "000000";
				when "101100010011" => data <= "000000";
				when "101100010100" => data <= "111111";
				when "101100010101" => data <= "100111";
				when "101100010110" => data <= "100111";
				when "101100010111" => data <= "111111";
				when "101100011000" => data <= "000000";
				when "101100011001" => data <= "000000";
				when "101100011010" => data <= "000000";
				when "101100011011" => data <= "000000";
				when "101100011100" => data <= "111111";
				when "101100011101" => data <= "100111";
				when "101100011110" => data <= "100111";
				when "101100011111" => data <= "111111";
				when "101100100000" => data <= "000000";
				when "101100100001" => data <= "000000";
				when "101100100010" => data <= "000000";
				when "101100100011" => data <= "000000";
				when "101100100100" => data <= "000000";
				when "101100100101" => data <= "000000";
				when "101100100110" => data <= "111111";
				when "101100100111" => data <= "100111";
				when "101100101000" => data <= "100111";
				when "101100101001" => data <= "100111";
				when "101100101010" => data <= "100111";
				when "101100101011" => data <= "100111";
				when "101100101100" => data <= "100111";
				when "101100101101" => data <= "100111";
				when "101100101110" => data <= "100111";
				when "101100101111" => data <= "100111";
				when "101100110000" => data <= "100111";
				when "101100110001" => data <= "111111";
				when "101100110010" => data <= "000000";
				when "101100110011" => data <= "000000";
				when "101100110100" => data <= "000000";
				when "101100110101" => data <= "000000";
				when "101100110110" => data <= "000000";
				when "101100110111" => data <= "000000";
				when "101100111000" => data <= "000000";
				when "101100111001" => data <= "000000";
				when "101100111010" => data <= "000000";
				when "101100111011" => data <= "000000";
				when "101100111100" => data <= "111111";
				when "101100111101" => data <= "100111";
				when "101100111110" => data <= "100111";
				when "101100111111" => data <= "111111";
				when "101101000000" => data <= "000000";
				when "101101000001" => data <= "000000";
				when "101101000010" => data <= "000000";
				when "101101000011" => data <= "000000";
				when "101101000100" => data <= "000000";
				when "101101000101" => data <= "000000";
				when "101101000110" => data <= "000000";
				when "101101000111" => data <= "000000";
				when "101101001000" => data <= "000000";
				when "101101001001" => data <= "000000";
				when "101101001010" => data <= "111111";
				when "101101001011" => data <= "100111";
				when "101101001100" => data <= "100111";
				when "101101001101" => data <= "111111";
				when "101101001110" => data <= "000000";
				when "101101001111" => data <= "000000";
				when "101101010000" => data <= "000000";
				when "101101010001" => data <= "000000";
				when "101101010010" => data <= "111111";
				when "101101010011" => data <= "100111";
				when "101101010100" => data <= "100111";
				when "101101010101" => data <= "111111";
				when "101101010110" => data <= "000000";
				when "101101010111" => data <= "000000";
				when "101101011000" => data <= "000000";
				when "101101011001" => data <= "000000";
				when "101101011010" => data <= "000000";
				when "101101011011" => data <= "000000";
				when "101101011100" => data <= "111111";
				when "101101011101" => data <= "100111";
				when "101101011110" => data <= "100111";
				when "101101011111" => data <= "100111";
				when "101101100000" => data <= "100111";
				when "101101100001" => data <= "100111";
				when "101101100010" => data <= "100111";
				when "101101100011" => data <= "100111";
				when "101101100100" => data <= "100111";
				when "101101100101" => data <= "100111";
				when "101101100110" => data <= "100111";
				when "101101100111" => data <= "111111";
				when "101101101000" => data <= "000000";
				when "101101101001" => data <= "000000";
				when "101101101010" => data <= "000000";
				when "101101101011" => data <= "000000";
				when "101101101100" => data <= "000000";
				when "101101101101" => data <= "000000";
				when "101101101110" => data <= "000000";
				when "101101101111" => data <= "000000";
				when "101101110000" => data <= "000000";
				when "101101110001" => data <= "000000";
				when "101101110010" => data <= "000000";
				when "101101110011" => data <= "000000";
				when "101101110100" => data <= "000000";
				when "101101110101" => data <= "000000";
				when "101101110110" => data <= "000000";
				when "101101110111" => data <= "000000";
				when "101101111000" => data <= "000000";
				when "101101111001" => data <= "000000";
				when "101101111010" => data <= "000000";
				when "101101111011" => data <= "000000";
				when "101101111100" => data <= "000000";
				when "101101111101" => data <= "000000";
				when "101101111110" => data <= "000000";
				when "101101111111" => data <= "000000";
				when "101110000000" => data <= "000000";
				when "101110000001" => data <= "000000";
				when "101110000010" => data <= "000000";
				when "101110000011" => data <= "000000";
				when "101110000100" => data <= "000000";
				when "101110000101" => data <= "000000";
				when "101110000110" => data <= "000000";
				when "101110000111" => data <= "000000";
				when "101110001000" => data <= "000000";
				when "101110001001" => data <= "000000";
				when "101110001010" => data <= "000000";
				when "101110001011" => data <= "000000";
				when "101110001100" => data <= "000000";
				when "101110001101" => data <= "000000";
				when "101110001110" => data <= "000000";
				when "101110001111" => data <= "000000";
				when "101110010000" => data <= "000000";
				when "101110010001" => data <= "000000";
				when "101110010010" => data <= "000000";
				when "101110010011" => data <= "000000";
				when "101110010100" => data <= "111111";
				when "101110010101" => data <= "100111";
				when "101110010110" => data <= "100111";
				when "101110010111" => data <= "111111";
				when "101110011000" => data <= "000000";
				when "101110011001" => data <= "000000";
				when "101110011010" => data <= "000000";
				when "101110011011" => data <= "000000";
				when "101110011100" => data <= "111111";
				when "101110011101" => data <= "100111";
				when "101110011110" => data <= "100111";
				when "101110011111" => data <= "111111";
				when "101110100000" => data <= "000000";
				when "101110100001" => data <= "000000";
				when "101110100010" => data <= "000000";
				when "101110100011" => data <= "000000";
				when "101110100100" => data <= "000000";
				when "101110100101" => data <= "000000";
				when "101110100110" => data <= "111111";
				when "101110100111" => data <= "100111";
				when "101110101000" => data <= "100111";
				when "101110101001" => data <= "100111";
				when "101110101010" => data <= "100111";
				when "101110101011" => data <= "100111";
				when "101110101100" => data <= "100111";
				when "101110101101" => data <= "100111";
				when "101110101110" => data <= "100111";
				when "101110101111" => data <= "100111";
				when "101110110000" => data <= "100111";
				when "101110110001" => data <= "111111";
				when "101110110010" => data <= "000000";
				when "101110110011" => data <= "000000";
				when "101110110100" => data <= "000000";
				when "101110110101" => data <= "000000";
				when "101110110110" => data <= "000000";
				when "101110110111" => data <= "000000";
				when "101110111000" => data <= "000000";
				when "101110111001" => data <= "000000";
				when "101110111010" => data <= "000000";
				when "101110111011" => data <= "000000";
				when "101110111100" => data <= "111111";
				when "101110111101" => data <= "100111";
				when "101110111110" => data <= "100111";
				when "101110111111" => data <= "111111";
				when "101111000000" => data <= "000000";
				when "101111000001" => data <= "000000";
				when "101111000010" => data <= "000000";
				when "101111000011" => data <= "000000";
				when "101111000100" => data <= "000000";
				when "101111000101" => data <= "000000";
				when "101111000110" => data <= "000000";
				when "101111000111" => data <= "000000";
				when "101111001000" => data <= "000000";
				when "101111001001" => data <= "000000";
				when "101111001010" => data <= "111111";
				when "101111001011" => data <= "100111";
				when "101111001100" => data <= "100111";
				when "101111001101" => data <= "111111";
				when "101111001110" => data <= "000000";
				when "101111001111" => data <= "000000";
				when "101111010000" => data <= "000000";
				when "101111010001" => data <= "000000";
				when "101111010010" => data <= "111111";
				when "101111010011" => data <= "100111";
				when "101111010100" => data <= "100111";
				when "101111010101" => data <= "111111";
				when "101111010110" => data <= "000000";
				when "101111010111" => data <= "000000";
				when "101111011000" => data <= "000000";
				when "101111011001" => data <= "000000";
				when "101111011010" => data <= "000000";
				when "101111011011" => data <= "000000";
				when "101111011100" => data <= "000000";
				when "101111011101" => data <= "111111";
				when "101111011110" => data <= "100111";
				when "101111011111" => data <= "100111";
				when "101111100000" => data <= "100111";
				when "101111100001" => data <= "100111";
				when "101111100010" => data <= "100111";
				when "101111100011" => data <= "100111";
				when "101111100100" => data <= "100111";
				when "101111100101" => data <= "100111";
				when "101111100110" => data <= "111111";
				when "101111100111" => data <= "000000";
				when "101111101000" => data <= "000000";
				when "101111101001" => data <= "000000";
				when "101111101010" => data <= "000000";
				when "101111101011" => data <= "000000";
				when "101111101100" => data <= "000000";
				when "101111101101" => data <= "000000";
				when "101111101110" => data <= "000000";
				when "101111101111" => data <= "000000";
				when "101111110000" => data <= "000000";
				when "101111110001" => data <= "000000";
				when "101111110010" => data <= "000000";
				when "101111110011" => data <= "000000";
				when "101111110100" => data <= "000000";
				when "101111110101" => data <= "000000";
				when "101111110110" => data <= "000000";
				when "101111110111" => data <= "000000";
				when "101111111000" => data <= "000000";
				when "101111111001" => data <= "000000";
				when "101111111010" => data <= "000000";
				when "101111111011" => data <= "000000";
				when "101111111100" => data <= "000000";
				when "101111111101" => data <= "000000";
				when "101111111110" => data <= "000000";
				when "101111111111" => data <= "000000";
				when "110000000000" => data <= "000000";
				when "110000000001" => data <= "000000";
				when "110000000010" => data <= "000000";
				when "110000000011" => data <= "000000";
				when "110000000100" => data <= "000000";
				when "110000000101" => data <= "000000";
				when "110000000110" => data <= "000000";
				when "110000000111" => data <= "000000";
				when "110000001000" => data <= "000000";
				when "110000001001" => data <= "000000";
				when "110000001010" => data <= "000000";
				when "110000001011" => data <= "000000";
				when "110000001100" => data <= "000000";
				when "110000001101" => data <= "000000";
				when "110000001110" => data <= "000000";
				when "110000001111" => data <= "000000";
				when "110000010000" => data <= "000000";
				when "110000010001" => data <= "000000";
				when "110000010010" => data <= "000000";
				when "110000010011" => data <= "000000";
				when "110000010100" => data <= "000000";
				when "110000010101" => data <= "111111";
				when "110000010110" => data <= "111111";
				when "110000010111" => data <= "000000";
				when "110000011000" => data <= "000000";
				when "110000011001" => data <= "000000";
				when "110000011010" => data <= "000000";
				when "110000011011" => data <= "000000";
				when "110000011100" => data <= "000000";
				when "110000011101" => data <= "111111";
				when "110000011110" => data <= "111111";
				when "110000011111" => data <= "000000";
				when "110000100000" => data <= "000000";
				when "110000100001" => data <= "000000";
				when "110000100010" => data <= "000000";
				when "110000100011" => data <= "000000";
				when "110000100100" => data <= "000000";
				when "110000100101" => data <= "000000";
				when "110000100110" => data <= "000000";
				when "110000100111" => data <= "111111";
				when "110000101000" => data <= "111111";
				when "110000101001" => data <= "111111";
				when "110000101010" => data <= "111111";
				when "110000101011" => data <= "111111";
				when "110000101100" => data <= "111111";
				when "110000101101" => data <= "111111";
				when "110000101110" => data <= "111111";
				when "110000101111" => data <= "111111";
				when "110000110000" => data <= "111111";
				when "110000110001" => data <= "000000";
				when "110000110010" => data <= "000000";
				when "110000110011" => data <= "000000";
				when "110000110100" => data <= "000000";
				when "110000110101" => data <= "000000";
				when "110000110110" => data <= "000000";
				when "110000110111" => data <= "000000";
				when "110000111000" => data <= "000000";
				when "110000111001" => data <= "000000";
				when "110000111010" => data <= "000000";
				when "110000111011" => data <= "000000";
				when "110000111100" => data <= "000000";
				when "110000111101" => data <= "111111";
				when "110000111110" => data <= "111111";
				when "110000111111" => data <= "000000";
				when "110001000000" => data <= "000000";
				when "110001000001" => data <= "000000";
				when "110001000010" => data <= "000000";
				when "110001000011" => data <= "000000";
				when "110001000100" => data <= "000000";
				when "110001000101" => data <= "000000";
				when "110001000110" => data <= "000000";
				when "110001000111" => data <= "000000";
				when "110001001000" => data <= "000000";
				when "110001001001" => data <= "000000";
				when "110001001010" => data <= "000000";
				when "110001001011" => data <= "111111";
				when "110001001100" => data <= "111111";
				when "110001001101" => data <= "000000";
				when "110001001110" => data <= "000000";
				when "110001001111" => data <= "000000";
				when "110001010000" => data <= "000000";
				when "110001010001" => data <= "000000";
				when "110001010010" => data <= "000000";
				when "110001010011" => data <= "111111";
				when "110001010100" => data <= "111111";
				when "110001010101" => data <= "000000";
				when "110001010110" => data <= "000000";
				when "110001010111" => data <= "000000";
				when "110001011000" => data <= "000000";
				when "110001011001" => data <= "000000";
				when "110001011010" => data <= "000000";
				when "110001011011" => data <= "000000";
				when "110001011100" => data <= "000000";
				when "110001011101" => data <= "000000";
				when "110001011110" => data <= "111111";
				when "110001011111" => data <= "111111";
				when "110001100000" => data <= "111111";
				when "110001100001" => data <= "111111";
				when "110001100010" => data <= "111111";
				when "110001100011" => data <= "111111";
				when "110001100100" => data <= "111111";
				when "110001100101" => data <= "111111";
				when "110001100110" => data <= "000000";
				when "110001100111" => data <= "000000";
				when "110001101000" => data <= "000000";
				when "110001101001" => data <= "000000";
				when "110001101010" => data <= "000000";
				when "110001101011" => data <= "000000";
				when "110001101100" => data <= "000000";
				when "110001101101" => data <= "000000";
				when "110001101110" => data <= "000000";
				when "110001101111" => data <= "000000";
				when "110001110000" => data <= "000000";
				when "110001110001" => data <= "000000";
				when "110001110010" => data <= "000000";
				when "110001110011" => data <= "000000";
				when "110001110100" => data <= "000000";
				when "110001110101" => data <= "000000";
				when "110001110110" => data <= "000000";
				when "110001110111" => data <= "000000";
				when "110001111000" => data <= "000000";
				when "110001111001" => data <= "000000";
				when "110001111010" => data <= "000000";
				when "110001111011" => data <= "000000";
				when "110001111100" => data <= "000000";
				when "110001111101" => data <= "000000";
				when "110001111110" => data <= "000000";
				when "110001111111" => data <= "000000";
				when "110010000000" => data <= "000000";
				when "110010000001" => data <= "000000";
				when "110010000010" => data <= "000000";
				when "110010000011" => data <= "000000";
				when "110010000100" => data <= "000000";
				when "110010000101" => data <= "000000";
				when "110010000110" => data <= "000000";
				when "110010000111" => data <= "000000";
				when "110010001000" => data <= "000000";
				when "110010001001" => data <= "000000";
				when "110010001010" => data <= "000000";
				when "110010001011" => data <= "000000";
				when "110010001100" => data <= "000000";
				when "110010001101" => data <= "000000";
				when "110010001110" => data <= "000000";
				when "110010001111" => data <= "000000";
				when "110010010000" => data <= "000000";
				when "110010010001" => data <= "000000";
				when "110010010010" => data <= "000000";
				when "110010010011" => data <= "000000";
				when "110010010100" => data <= "000000";
				when "110010010101" => data <= "000000";
				when "110010010110" => data <= "000000";
				when "110010010111" => data <= "000000";
				when "110010011000" => data <= "000000";
				when "110010011001" => data <= "000000";
				when "110010011010" => data <= "000000";
				when "110010011011" => data <= "000000";
				when "110010011100" => data <= "000000";
				when "110010011101" => data <= "000000";
				when "110010011110" => data <= "000000";
				when "110010011111" => data <= "000000";
				when "110010100000" => data <= "000000";
				when "110010100001" => data <= "000000";
				when "110010100010" => data <= "000000";
				when "110010100011" => data <= "000000";
				when "110010100100" => data <= "000000";
				when "110010100101" => data <= "000000";
				when "110010100110" => data <= "000000";
				when "110010100111" => data <= "000000";
				when "110010101000" => data <= "000000";
				when "110010101001" => data <= "000000";
				when "110010101010" => data <= "000000";
				when "110010101011" => data <= "000000";
				when "110010101100" => data <= "000000";
				when "110010101101" => data <= "000000";
				when "110010101110" => data <= "000000";
				when "110010101111" => data <= "000000";
				when "110010110000" => data <= "000000";
				when "110010110001" => data <= "000000";
				when "110010110010" => data <= "000000";
				when "110010110011" => data <= "000000";
				when "110010110100" => data <= "000000";
				when "110010110101" => data <= "000000";
				when "110010110110" => data <= "000000";
				when "110010110111" => data <= "000000";
				when "110010111000" => data <= "000000";
				when "110010111001" => data <= "000000";
				when "110010111010" => data <= "000000";
				when "110010111011" => data <= "000000";
				when "110010111100" => data <= "000000";
				when "110010111101" => data <= "000000";
				when "110010111110" => data <= "000000";
				when "110010111111" => data <= "000000";
				when "110011000000" => data <= "000000";
				when "110011000001" => data <= "000000";
				when "110011000010" => data <= "000000";
				when "110011000011" => data <= "000000";
				when "110011000100" => data <= "000000";
				when "110011000101" => data <= "000000";
				when "110011000110" => data <= "000000";
				when "110011000111" => data <= "000000";
				when "110011001000" => data <= "000000";
				when "110011001001" => data <= "000000";
				when "110011001010" => data <= "000000";
				when "110011001011" => data <= "000000";
				when "110011001100" => data <= "000000";
				when "110011001101" => data <= "000000";
				when "110011001110" => data <= "000000";
				when "110011001111" => data <= "000000";
				when "110011010000" => data <= "000000";
				when "110011010001" => data <= "000000";
				when "110011010010" => data <= "000000";
				when "110011010011" => data <= "000000";
				when "110011010100" => data <= "000000";
				when "110011010101" => data <= "000000";
				when "110011010110" => data <= "000000";
				when "110011010111" => data <= "000000";
				when "110011011000" => data <= "000000";
				when "110011011001" => data <= "000000";
				when "110011011010" => data <= "000000";
				when "110011011011" => data <= "000000";
				when "110011011100" => data <= "000000";
				when "110011011101" => data <= "000000";
				when "110011011110" => data <= "000000";
				when "110011011111" => data <= "000000";
				when "110011100000" => data <= "000000";
				when "110011100001" => data <= "000000";
				when "110011100010" => data <= "000000";
				when "110011100011" => data <= "000000";
				when "110011100100" => data <= "000000";
				when "110011100101" => data <= "000000";
				when "110011100110" => data <= "000000";
				when "110011100111" => data <= "000000";
				when "110011101000" => data <= "000000";
				when "110011101001" => data <= "000000";
				when "110011101010" => data <= "000000";
				when "110011101011" => data <= "000000";
				when "110011101100" => data <= "000000";
				when "110011101101" => data <= "000000";
				when "110011101110" => data <= "000000";
				when "110011101111" => data <= "000000";
				when "110011110000" => data <= "000000";
				when "110011110001" => data <= "000000";
				when "110011110010" => data <= "000000";
				when "110011110011" => data <= "000000";
				when "110011110100" => data <= "000000";
				when "110011110101" => data <= "000000";
				when "110011110110" => data <= "000000";
				when "110011110111" => data <= "000000";
				when "110011111000" => data <= "000000";
				when "110011111001" => data <= "000000";
				when "110011111010" => data <= "000000";
				when "110011111011" => data <= "000000";
				when "110011111100" => data <= "000000";
				when "110011111101" => data <= "000000";
				when "110011111110" => data <= "000000";
				when "110011111111" => data <= "000000";
				when "110100000000" => data <= "000000";
				when "110100000001" => data <= "000000";
				when "110100000010" => data <= "000000";
				when "110100000011" => data <= "000000";
				when "110100000100" => data <= "000000";
				when "110100000101" => data <= "000000";
				when "110100000110" => data <= "000000";
				when "110100000111" => data <= "000000";
				when "110100001000" => data <= "000000";
				when "110100001001" => data <= "000000";
				when "110100001010" => data <= "000000";
				when "110100001011" => data <= "000000";
				when "110100001100" => data <= "000000";
				when "110100001101" => data <= "000000";
				when "110100001110" => data <= "000000";
				when "110100001111" => data <= "000000";
				when "110100010000" => data <= "000000";
				when "110100010001" => data <= "000000";
				when "110100010010" => data <= "000000";
				when "110100010011" => data <= "000000";
				when "110100010100" => data <= "000000";
				when "110100010101" => data <= "000000";
				when "110100010110" => data <= "000000";
				when "110100010111" => data <= "000000";
				when "110100011000" => data <= "000000";
				when "110100011001" => data <= "000000";
				when "110100011010" => data <= "000000";
				when "110100011011" => data <= "000000";
				when "110100011100" => data <= "000000";
				when "110100011101" => data <= "000000";
				when "110100011110" => data <= "000000";
				when "110100011111" => data <= "000000";
				when "110100100000" => data <= "000000";
				when "110100100001" => data <= "000000";
				when "110100100010" => data <= "000000";
				when "110100100011" => data <= "000000";
				when "110100100100" => data <= "000000";
				when "110100100101" => data <= "000000";
				when "110100100110" => data <= "000000";
				when "110100100111" => data <= "000000";
				when "110100101000" => data <= "000000";
				when "110100101001" => data <= "000000";
				when "110100101010" => data <= "000000";
				when "110100101011" => data <= "000000";
				when "110100101100" => data <= "000000";
				when "110100101101" => data <= "000000";
				when "110100101110" => data <= "000000";
				when "110100101111" => data <= "000000";
				when "110100110000" => data <= "000000";
				when "110100110001" => data <= "000000";
				when "110100110010" => data <= "000000";
				when "110100110011" => data <= "000000";
				when "110100110100" => data <= "000000";
				when "110100110101" => data <= "000000";
				when "110100110110" => data <= "000000";
				when "110100110111" => data <= "000000";
				when "110100111000" => data <= "000000";
				when "110100111001" => data <= "000000";
				when "110100111010" => data <= "000000";
				when "110100111011" => data <= "000000";
				when "110100111100" => data <= "000000";
				when "110100111101" => data <= "000000";
				when "110100111110" => data <= "000000";
				when "110100111111" => data <= "000000";
				when "110101000000" => data <= "000000";
				when "110101000001" => data <= "000000";
				when "110101000010" => data <= "000000";
				when "110101000011" => data <= "000000";
				when "110101000100" => data <= "000000";
				when "110101000101" => data <= "000000";
				when "110101000110" => data <= "000000";
				when "110101000111" => data <= "000000";
				when "110101001000" => data <= "000000";
				when "110101001001" => data <= "000000";
				when "110101001010" => data <= "000000";
				when "110101001011" => data <= "000000";
				when "110101001100" => data <= "000000";
				when "110101001101" => data <= "000000";
				when "110101001110" => data <= "000000";
				when "110101001111" => data <= "000000";
				when "110101010000" => data <= "000000";
				when "110101010001" => data <= "000000";
				when "110101010010" => data <= "000000";
				when "110101010011" => data <= "000000";
				when "110101010100" => data <= "000000";
				when "110101010101" => data <= "000000";
				when "110101010110" => data <= "000000";
				when "110101010111" => data <= "000000";
				when "110101011000" => data <= "000000";
				when "110101011001" => data <= "000000";
				when "110101011010" => data <= "000000";
				when "110101011011" => data <= "000000";
				when "110101011100" => data <= "000000";
				when "110101011101" => data <= "000000";
				when "110101011110" => data <= "000000";
				when "110101011111" => data <= "000000";
				when "110101100000" => data <= "000000";
				when "110101100001" => data <= "000000";
				when "110101100010" => data <= "000000";
				when "110101100011" => data <= "000000";
				when "110101100100" => data <= "000000";
				when "110101100101" => data <= "000000";
				when "110101100110" => data <= "000000";
				when "110101100111" => data <= "000000";
				when "110101101000" => data <= "000000";
				when "110101101001" => data <= "000000";
				when "110101101010" => data <= "000000";
				when "110101101011" => data <= "000000";
				when "110101101100" => data <= "000000";
				when "110101101101" => data <= "000000";
				when "110101101110" => data <= "000000";
				when "110101101111" => data <= "000000";
				when "110101110000" => data <= "000000";
				when "110101110001" => data <= "000000";
				when "110101110010" => data <= "000000";
				when "110101110011" => data <= "000000";
				when "110101110100" => data <= "000000";
				when "110101110101" => data <= "000000";
				when "110101110110" => data <= "000000";
				when "110101110111" => data <= "000000";
				when "110101111000" => data <= "000000";
				when "110101111001" => data <= "000000";
				when "110101111010" => data <= "000000";
				when "110101111011" => data <= "000000";
				when "110101111100" => data <= "000000";
				when "110101111101" => data <= "000000";
				when "110101111110" => data <= "000000";
				when "110101111111" => data <= "000000";
				when "110110000000" => data <= "000000";
				when "110110000001" => data <= "000000";
				when "110110000010" => data <= "000000";
				when "110110000011" => data <= "000000";
				when "110110000100" => data <= "000000";
				when "110110000101" => data <= "000000";
				when "110110000110" => data <= "000000";
				when "110110000111" => data <= "000000";
				when "110110001000" => data <= "000000";
				when "110110001001" => data <= "000000";
				when "110110001010" => data <= "000000";
				when "110110001011" => data <= "000000";
				when "110110001100" => data <= "000000";
				when "110110001101" => data <= "000000";
				when "110110001110" => data <= "000000";
				when "110110001111" => data <= "000000";
				when "110110010000" => data <= "000000";
				when "110110010001" => data <= "000000";
				when "110110010010" => data <= "000000";
				when "110110010011" => data <= "000000";
				when "110110010100" => data <= "000000";
				when "110110010101" => data <= "000000";
				when "110110010110" => data <= "000000";
				when "110110010111" => data <= "000000";
				when "110110011000" => data <= "000000";
				when "110110011001" => data <= "000000";
				when "110110011010" => data <= "000000";
				when "110110011011" => data <= "000000";
				when "110110011100" => data <= "000000";
				when "110110011101" => data <= "000000";
				when "110110011110" => data <= "000000";
				when "110110011111" => data <= "000000";
				when "110110100000" => data <= "000000";
				when "110110100001" => data <= "000000";
				when "110110100010" => data <= "000000";
				when "110110100011" => data <= "000000";
				when "110110100100" => data <= "000000";
				when "110110100101" => data <= "000000";
				when "110110100110" => data <= "000000";
				when "110110100111" => data <= "000000";
				when "110110101000" => data <= "000000";
				when "110110101001" => data <= "000000";
				when "110110101010" => data <= "000000";
				when "110110101011" => data <= "000000";
				when "110110101100" => data <= "000000";
				when "110110101101" => data <= "000000";
				when "110110101110" => data <= "000000";
				when "110110101111" => data <= "000000";
				when "110110110000" => data <= "000000";
				when "110110110001" => data <= "000000";
				when "110110110010" => data <= "000000";
				when "110110110011" => data <= "000000";
				when "110110110100" => data <= "000000";
				when "110110110101" => data <= "000000";
				when "110110110110" => data <= "000000";
				when "110110110111" => data <= "000000";
				when "110110111000" => data <= "000000";
				when "110110111001" => data <= "000000";
				when "110110111010" => data <= "000000";
				when "110110111011" => data <= "000000";
				when "110110111100" => data <= "000000";
				when "110110111101" => data <= "000000";
				when "110110111110" => data <= "000000";
				when "110110111111" => data <= "000000";
				when "110111000000" => data <= "000000";
				when "110111000001" => data <= "000000";
				when "110111000010" => data <= "000000";
				when "110111000011" => data <= "000000";
				when "110111000100" => data <= "000000";
				when "110111000101" => data <= "000000";
				when "110111000110" => data <= "000000";
				when "110111000111" => data <= "000000";
				when "110111001000" => data <= "000000";
				when "110111001001" => data <= "000000";
				when "110111001010" => data <= "000000";
				when "110111001011" => data <= "000000";
				when "110111001100" => data <= "000000";
				when "110111001101" => data <= "000000";
				when "110111001110" => data <= "000000";
				when "110111001111" => data <= "000000";
				when "110111010000" => data <= "000000";
				when "110111010001" => data <= "000000";
				when "110111010010" => data <= "000000";
				when "110111010011" => data <= "000000";
				when "110111010100" => data <= "000000";
				when "110111010101" => data <= "000000";
				when "110111010110" => data <= "000000";
				when "110111010111" => data <= "000000";
				when "110111011000" => data <= "000000";
				when "110111011001" => data <= "000000";
				when "110111011010" => data <= "000000";
				when "110111011011" => data <= "000000";
				when "110111011100" => data <= "000000";
				when "110111011101" => data <= "000000";
				when "110111011110" => data <= "000000";
				when "110111011111" => data <= "000000";
				when "110111100000" => data <= "000000";
				when "110111100001" => data <= "000000";
				when "110111100010" => data <= "000000";
				when "110111100011" => data <= "000000";
				when "110111100100" => data <= "000000";
				when "110111100101" => data <= "000000";
				when "110111100110" => data <= "000000";
				when "110111100111" => data <= "000000";
				when "110111101000" => data <= "000000";
				when "110111101001" => data <= "000000";
				when "110111101010" => data <= "000000";
				when "110111101011" => data <= "000000";
				when "110111101100" => data <= "000000";
				when "110111101101" => data <= "000000";
				when "110111101110" => data <= "000000";
				when "110111101111" => data <= "000000";
				when "110111110000" => data <= "000000";
				when "110111110001" => data <= "000000";
				when "110111110010" => data <= "000000";
				when "110111110011" => data <= "000000";
				when "110111110100" => data <= "000000";
				when "110111110101" => data <= "000000";
				when "110111110110" => data <= "000000";
				when "110111110111" => data <= "000000";
				when "110111111000" => data <= "000000";
				when "110111111001" => data <= "000000";
				when "110111111010" => data <= "000000";
				when "110111111011" => data <= "000000";
				when "110111111100" => data <= "000000";
				when "110111111101" => data <= "000000";
				when "110111111110" => data <= "000000";
				when "110111111111" => data <= "000000";
				when "111000000000" => data <= "000000";
				when "111000000001" => data <= "000000";
				when "111000000010" => data <= "000000";
				when "111000000011" => data <= "000000";
				when "111000000100" => data <= "000000";
				when "111000000101" => data <= "000000";
				when "111000000110" => data <= "000000";
				when "111000000111" => data <= "000000";
				when "111000001000" => data <= "000000";
				when "111000001001" => data <= "000000";
				when "111000001010" => data <= "000000";
				when "111000001011" => data <= "000000";
				when "111000001100" => data <= "000000";
				when "111000001101" => data <= "000000";
				when "111000001110" => data <= "000000";
				when "111000001111" => data <= "000000";
				when "111000010000" => data <= "000000";
				when "111000010001" => data <= "000000";
				when "111000010010" => data <= "000000";
				when "111000010011" => data <= "000000";
				when "111000010100" => data <= "000000";
				when "111000010101" => data <= "000000";
				when "111000010110" => data <= "000000";
				when "111000010111" => data <= "000000";
				when "111000011000" => data <= "000000";
				when "111000011001" => data <= "000000";
				when "111000011010" => data <= "000000";
				when "111000011011" => data <= "000000";
				when "111000011100" => data <= "000000";
				when "111000011101" => data <= "000000";
				when "111000011110" => data <= "000000";
				when "111000011111" => data <= "000000";
				when "111000100000" => data <= "000000";
				when "111000100001" => data <= "000000";
				when "111000100010" => data <= "000000";
				when "111000100011" => data <= "000000";
				when "111000100100" => data <= "000000";
				when "111000100101" => data <= "000000";
				when "111000100110" => data <= "000000";
				when "111000100111" => data <= "000000";
				when "111000101000" => data <= "000000";
				when "111000101001" => data <= "000000";
				when "111000101010" => data <= "000000";
				when "111000101011" => data <= "000000";
				when "111000101100" => data <= "000000";
				when "111000101101" => data <= "000000";
				when "111000101110" => data <= "000000";
				when "111000101111" => data <= "000000";
				when "111000110000" => data <= "000000";
				when "111000110001" => data <= "000000";
				when "111000110010" => data <= "000000";
				when "111000110011" => data <= "000000";
				when "111000110100" => data <= "000000";
				when "111000110101" => data <= "000000";
				when "111000110110" => data <= "000000";
				when "111000110111" => data <= "000000";
				when "111000111000" => data <= "000000";
				when "111000111001" => data <= "000000";
				when "111000111010" => data <= "000000";
				when "111000111011" => data <= "000000";
				when "111000111100" => data <= "000000";
				when "111000111101" => data <= "000000";
				when "111000111110" => data <= "000000";
				when "111000111111" => data <= "000000";
				when "111001000000" => data <= "000000";
				when "111001000001" => data <= "000000";
				when "111001000010" => data <= "000000";
				when "111001000011" => data <= "000000";
				when "111001000100" => data <= "000000";
				when "111001000101" => data <= "000000";
				when "111001000110" => data <= "000000";
				when "111001000111" => data <= "000000";
				when "111001001000" => data <= "000000";
				when "111001001001" => data <= "000000";
				when "111001001010" => data <= "000000";
				when "111001001011" => data <= "000000";
				when "111001001100" => data <= "000000";
				when "111001001101" => data <= "000000";
				when "111001001110" => data <= "000000";
				when "111001001111" => data <= "000000";
				when "111001010000" => data <= "000000";
				when "111001010001" => data <= "000000";
				when "111001010010" => data <= "000000";
				when "111001010011" => data <= "000000";
				when "111001010100" => data <= "000000";
				when "111001010101" => data <= "000000";
				when "111001010110" => data <= "000000";
				when "111001010111" => data <= "000000";
				when "111001011000" => data <= "000000";
				when "111001011001" => data <= "000000";
				when "111001011010" => data <= "000000";
				when "111001011011" => data <= "000000";
				when "111001011100" => data <= "000000";
				when "111001011101" => data <= "000000";
				when "111001011110" => data <= "000000";
				when "111001011111" => data <= "000000";
				when "111001100000" => data <= "000000";
				when "111001100001" => data <= "000000";
				when "111001100010" => data <= "000000";
				when "111001100011" => data <= "000000";
				when "111001100100" => data <= "000000";
				when "111001100101" => data <= "000000";
				when "111001100110" => data <= "000000";
				when "111001100111" => data <= "000000";
				when "111001101000" => data <= "000000";
				when "111001101001" => data <= "000000";
				when "111001101010" => data <= "000000";
				when "111001101011" => data <= "000000";
				when "111001101100" => data <= "000000";
				when "111001101101" => data <= "000000";
				when "111001101110" => data <= "000000";
				when "111001101111" => data <= "000000";
				when "111001110000" => data <= "000000";
				when "111001110001" => data <= "000000";
				when "111001110010" => data <= "000000";
				when "111001110011" => data <= "000000";
				when "111001110100" => data <= "000000";
				when "111001110101" => data <= "000000";
				when "111001110110" => data <= "000000";
				when "111001110111" => data <= "000000";
				when "111001111000" => data <= "000000";
				when "111001111001" => data <= "000000";
				when "111001111010" => data <= "000000";
				when "111001111011" => data <= "000000";
				when "111001111100" => data <= "000000";
				when "111001111101" => data <= "000000";
				when "111001111110" => data <= "000000";
				when "111001111111" => data <= "000000";
				when "111010000000" => data <= "000000";
				when "111010000001" => data <= "000000";
				when "111010000010" => data <= "000000";
				when "111010000011" => data <= "000000";
				when "111010000100" => data <= "000000";
				when "111010000101" => data <= "000000";
				when "111010000110" => data <= "000000";
				when "111010000111" => data <= "000000";
				when "111010001000" => data <= "000000";
				when "111010001001" => data <= "000000";
				when "111010001010" => data <= "000000";
				when "111010001011" => data <= "000000";
				when "111010001100" => data <= "000000";
				when "111010001101" => data <= "000000";
				when "111010001110" => data <= "111111";
				when "111010001111" => data <= "111111";
				when "111010010000" => data <= "111111";
				when "111010010001" => data <= "111111";
				when "111010010010" => data <= "111111";
				when "111010010011" => data <= "111111";
				when "111010010100" => data <= "111111";
				when "111010010101" => data <= "111111";
				when "111010010110" => data <= "000000";
				when "111010010111" => data <= "000000";
				when "111010011000" => data <= "000000";
				when "111010011001" => data <= "000000";
				when "111010011010" => data <= "000000";
				when "111010011011" => data <= "000000";
				when "111010011100" => data <= "000000";
				when "111010011101" => data <= "000000";
				when "111010011110" => data <= "000000";
				when "111010011111" => data <= "111111";
				when "111010100000" => data <= "111111";
				when "111010100001" => data <= "000000";
				when "111010100010" => data <= "000000";
				when "111010100011" => data <= "000000";
				when "111010100100" => data <= "000000";
				when "111010100101" => data <= "000000";
				when "111010100110" => data <= "000000";
				when "111010100111" => data <= "111111";
				when "111010101000" => data <= "111111";
				when "111010101001" => data <= "000000";
				when "111010101010" => data <= "000000";
				when "111010101011" => data <= "000000";
				when "111010101100" => data <= "000000";
				when "111010101101" => data <= "000000";
				when "111010101110" => data <= "000000";
				when "111010101111" => data <= "111111";
				when "111010110000" => data <= "111111";
				when "111010110001" => data <= "111111";
				when "111010110010" => data <= "111111";
				when "111010110011" => data <= "111111";
				when "111010110100" => data <= "111111";
				when "111010110101" => data <= "111111";
				when "111010110110" => data <= "111111";
				when "111010110111" => data <= "111111";
				when "111010111000" => data <= "111111";
				when "111010111001" => data <= "111111";
				when "111010111010" => data <= "111111";
				when "111010111011" => data <= "000000";
				when "111010111100" => data <= "000000";
				when "111010111101" => data <= "000000";
				when "111010111110" => data <= "000000";
				when "111010111111" => data <= "000000";
				when "111011000000" => data <= "111111";
				when "111011000001" => data <= "111111";
				when "111011000010" => data <= "000000";
				when "111011000011" => data <= "000000";
				when "111011000100" => data <= "000000";
				when "111011000101" => data <= "000000";
				when "111011000110" => data <= "000000";
				when "111011000111" => data <= "000000";
				when "111011001000" => data <= "111111";
				when "111011001001" => data <= "111111";
				when "111011001010" => data <= "000000";
				when "111011001011" => data <= "000000";
				when "111011001100" => data <= "000000";
				when "111011001101" => data <= "000000";
				when "111011001110" => data <= "000000";
				when "111011001111" => data <= "000000";
				when "111011010000" => data <= "111111";
				when "111011010001" => data <= "111111";
				when "111011010010" => data <= "000000";
				when "111011010011" => data <= "000000";
				when "111011010100" => data <= "000000";
				when "111011010101" => data <= "000000";
				when "111011010110" => data <= "000000";
				when "111011010111" => data <= "000000";
				when "111011011000" => data <= "111111";
				when "111011011001" => data <= "111111";
				when "111011011010" => data <= "000000";
				when "111011011011" => data <= "000000";
				when "111011011100" => data <= "000000";
				when "111011011101" => data <= "000000";
				when "111011011110" => data <= "000000";
				when "111011011111" => data <= "000000";
				when "111011100000" => data <= "000000";
				when "111011100001" => data <= "000000";
				when "111011100010" => data <= "111111";
				when "111011100011" => data <= "111111";
				when "111011100100" => data <= "000000";
				when "111011100101" => data <= "000000";
				when "111011100110" => data <= "000000";
				when "111011100111" => data <= "000000";
				when "111011101000" => data <= "000000";
				when "111011101001" => data <= "000000";
				when "111011101010" => data <= "111111";
				when "111011101011" => data <= "111111";
				when "111011101100" => data <= "000000";
				when "111011101101" => data <= "000000";
				when "111011101110" => data <= "000000";
				when "111011101111" => data <= "000000";
				when "111011110000" => data <= "000000";
				when "111011110001" => data <= "000000";
				when "111011110010" => data <= "000000";
				when "111011110011" => data <= "000000";
				when "111011110100" => data <= "000000";
				when "111011110101" => data <= "000000";
				when "111011110110" => data <= "000000";
				when "111011110111" => data <= "000000";
				when "111011111000" => data <= "000000";
				when "111011111001" => data <= "000000";
				when "111011111010" => data <= "000000";
				when "111011111011" => data <= "000000";
				when "111011111100" => data <= "000000";
				when "111011111101" => data <= "000000";
				when "111011111110" => data <= "000000";
				when "111011111111" => data <= "000000";
				when "111100000000" => data <= "000000";
				when "111100000001" => data <= "000000";
				when "111100000010" => data <= "000000";
				when "111100000011" => data <= "000000";
				when "111100000100" => data <= "000000";
				when "111100000101" => data <= "000000";
				when "111100000110" => data <= "000000";
				when "111100000111" => data <= "000000";
				when "111100001000" => data <= "000000";
				when "111100001001" => data <= "000000";
				when "111100001010" => data <= "000000";
				when "111100001011" => data <= "000000";
				when "111100001100" => data <= "000000";
				when "111100001101" => data <= "111111";
				when "111100001110" => data <= "010010";
				when "111100001111" => data <= "010010";
				when "111100010000" => data <= "010010";
				when "111100010001" => data <= "010010";
				when "111100010010" => data <= "010010";
				when "111100010011" => data <= "010010";
				when "111100010100" => data <= "010010";
				when "111100010101" => data <= "010010";
				when "111100010110" => data <= "111111";
				when "111100010111" => data <= "000000";
				when "111100011000" => data <= "000000";
				when "111100011001" => data <= "000000";
				when "111100011010" => data <= "000000";
				when "111100011011" => data <= "000000";
				when "111100011100" => data <= "000000";
				when "111100011101" => data <= "000000";
				when "111100011110" => data <= "111111";
				when "111100011111" => data <= "010010";
				when "111100100000" => data <= "010010";
				when "111100100001" => data <= "111111";
				when "111100100010" => data <= "000000";
				when "111100100011" => data <= "000000";
				when "111100100100" => data <= "000000";
				when "111100100101" => data <= "000000";
				when "111100100110" => data <= "111111";
				when "111100100111" => data <= "010010";
				when "111100101000" => data <= "010010";
				when "111100101001" => data <= "111111";
				when "111100101010" => data <= "000000";
				when "111100101011" => data <= "000000";
				when "111100101100" => data <= "000000";
				when "111100101101" => data <= "000000";
				when "111100101110" => data <= "111111";
				when "111100101111" => data <= "010010";
				when "111100110000" => data <= "010010";
				when "111100110001" => data <= "010010";
				when "111100110010" => data <= "010010";
				when "111100110011" => data <= "010010";
				when "111100110100" => data <= "010010";
				when "111100110101" => data <= "010010";
				when "111100110110" => data <= "010010";
				when "111100110111" => data <= "010010";
				when "111100111000" => data <= "010010";
				when "111100111001" => data <= "010010";
				when "111100111010" => data <= "010010";
				when "111100111011" => data <= "111111";
				when "111100111100" => data <= "000000";
				when "111100111101" => data <= "000000";
				when "111100111110" => data <= "000000";
				when "111100111111" => data <= "111111";
				when "111101000000" => data <= "010010";
				when "111101000001" => data <= "010010";
				when "111101000010" => data <= "111111";
				when "111101000011" => data <= "000000";
				when "111101000100" => data <= "000000";
				when "111101000101" => data <= "000000";
				when "111101000110" => data <= "000000";
				when "111101000111" => data <= "111111";
				when "111101001000" => data <= "010010";
				when "111101001001" => data <= "010010";
				when "111101001010" => data <= "111111";
				when "111101001011" => data <= "000000";
				when "111101001100" => data <= "000000";
				when "111101001101" => data <= "000000";
				when "111101001110" => data <= "000000";
				when "111101001111" => data <= "111111";
				when "111101010000" => data <= "010010";
				when "111101010001" => data <= "010010";
				when "111101010010" => data <= "111111";
				when "111101010011" => data <= "000000";
				when "111101010100" => data <= "000000";
				when "111101010101" => data <= "000000";
				when "111101010110" => data <= "000000";
				when "111101010111" => data <= "111111";
				when "111101011000" => data <= "010010";
				when "111101011001" => data <= "010010";
				when "111101011010" => data <= "111111";
				when "111101011011" => data <= "000000";
				when "111101011100" => data <= "000000";
				when "111101011101" => data <= "000000";
				when "111101011110" => data <= "000000";
				when "111101011111" => data <= "000000";
				when "111101100000" => data <= "000000";
				when "111101100001" => data <= "111111";
				when "111101100010" => data <= "010010";
				when "111101100011" => data <= "010010";
				when "111101100100" => data <= "111111";
				when "111101100101" => data <= "000000";
				when "111101100110" => data <= "000000";
				when "111101100111" => data <= "000000";
				when "111101101000" => data <= "000000";
				when "111101101001" => data <= "111111";
				when "111101101010" => data <= "010010";
				when "111101101011" => data <= "010010";
				when "111101101100" => data <= "111111";
				when "111101101101" => data <= "000000";
				when "111101101110" => data <= "000000";
				when "111101101111" => data <= "000000";
				when "111101110000" => data <= "000000";
				when "111101110001" => data <= "000000";
				when "111101110010" => data <= "000000";
				when "111101110011" => data <= "000000";
				when "111101110100" => data <= "000000";
				when "111101110101" => data <= "000000";
				when "111101110110" => data <= "000000";
				when "111101110111" => data <= "000000";
				when "111101111000" => data <= "000000";
				when "111101111001" => data <= "000000";
				when "111101111010" => data <= "000000";
				when "111101111011" => data <= "000000";
				when "111101111100" => data <= "000000";
				when "111101111101" => data <= "000000";
				when "111101111110" => data <= "000000";
				when "111101111111" => data <= "000000";
				when "111110000000" => data <= "000000";
				when "111110000001" => data <= "000000";
				when "111110000010" => data <= "000000";
				when "111110000011" => data <= "000000";
				when "111110000100" => data <= "000000";
				when "111110000101" => data <= "000000";
				when "111110000110" => data <= "000000";
				when "111110000111" => data <= "000000";
				when "111110001000" => data <= "000000";
				when "111110001001" => data <= "000000";
				when "111110001010" => data <= "000000";
				when "111110001011" => data <= "000000";
				when "111110001100" => data <= "000000";
				when "111110001101" => data <= "111111";
				when "111110001110" => data <= "010010";
				when "111110001111" => data <= "010010";
				when "111110010000" => data <= "010010";
				when "111110010001" => data <= "010010";
				when "111110010010" => data <= "010010";
				when "111110010011" => data <= "010010";
				when "111110010100" => data <= "010010";
				when "111110010101" => data <= "010010";
				when "111110010110" => data <= "111111";
				when "111110010111" => data <= "111111";
				when "111110011000" => data <= "000000";
				when "111110011001" => data <= "000000";
				when "111110011010" => data <= "000000";
				when "111110011011" => data <= "000000";
				when "111110011100" => data <= "000000";
				when "111110011101" => data <= "000000";
				when "111110011110" => data <= "111111";
				when "111110011111" => data <= "010010";
				when "111110100000" => data <= "010010";
				when "111110100001" => data <= "111111";
				when "111110100010" => data <= "000000";
				when "111110100011" => data <= "000000";
				when "111110100100" => data <= "000000";
				when "111110100101" => data <= "000000";
				when "111110100110" => data <= "111111";
				when "111110100111" => data <= "010010";
				when "111110101000" => data <= "010010";
				when "111110101001" => data <= "111111";
				when "111110101010" => data <= "000000";
				when "111110101011" => data <= "000000";
				when "111110101100" => data <= "000000";
				when "111110101101" => data <= "000000";
				when "111110101110" => data <= "111111";
				when "111110101111" => data <= "010010";
				when "111110110000" => data <= "010010";
				when "111110110001" => data <= "010010";
				when "111110110010" => data <= "010010";
				when "111110110011" => data <= "010010";
				when "111110110100" => data <= "010010";
				when "111110110101" => data <= "010010";
				when "111110110110" => data <= "010010";
				when "111110110111" => data <= "010010";
				when "111110111000" => data <= "010010";
				when "111110111001" => data <= "010010";
				when "111110111010" => data <= "010010";
				when "111110111011" => data <= "111111";
				when "111110111100" => data <= "000000";
				when "111110111101" => data <= "000000";
				when "111110111110" => data <= "000000";
				when "111110111111" => data <= "111111";
				when "111111000000" => data <= "010010";
				when "111111000001" => data <= "010010";
				when "111111000010" => data <= "111111";
				when "111111000011" => data <= "000000";
				when "111111000100" => data <= "000000";
				when "111111000101" => data <= "000000";
				when "111111000110" => data <= "000000";
				when "111111000111" => data <= "111111";
				when "111111001000" => data <= "010010";
				when "111111001001" => data <= "010010";
				when "111111001010" => data <= "111111";
				when "111111001011" => data <= "000000";
				when "111111001100" => data <= "000000";
				when "111111001101" => data <= "000000";
				when "111111001110" => data <= "000000";
				when "111111001111" => data <= "111111";
				when "111111010000" => data <= "010010";
				when "111111010001" => data <= "010010";
				when "111111010010" => data <= "111111";
				when "111111010011" => data <= "000000";
				when "111111010100" => data <= "000000";
				when "111111010101" => data <= "000000";
				when "111111010110" => data <= "000000";
				when "111111010111" => data <= "111111";
				when "111111011000" => data <= "010010";
				when "111111011001" => data <= "010010";
				when "111111011010" => data <= "111111";
				when "111111011011" => data <= "000000";
				when "111111011100" => data <= "000000";
				when "111111011101" => data <= "000000";
				when "111111011110" => data <= "000000";
				when "111111011111" => data <= "000000";
				when "111111100000" => data <= "000000";
				when "111111100001" => data <= "111111";
				when "111111100010" => data <= "010010";
				when "111111100011" => data <= "010010";
				when "111111100100" => data <= "111111";
				when "111111100101" => data <= "111111";
				when "111111100110" => data <= "000000";
				when "111111100111" => data <= "000000";
				when "111111101000" => data <= "111111";
				when "111111101001" => data <= "111111";
				when "111111101010" => data <= "010010";
				when "111111101011" => data <= "010010";
				when "111111101100" => data <= "111111";
				when "111111101101" => data <= "000000";
				when "111111101110" => data <= "000000";
				when "111111101111" => data <= "000000";
				when "111111110000" => data <= "000000";
				when "111111110001" => data <= "000000";
				when "111111110010" => data <= "000000";
				when "111111110011" => data <= "000000";
				when "111111110100" => data <= "000000";
				when "111111110101" => data <= "000000";
				when "111111110110" => data <= "000000";
				when "111111110111" => data <= "000000";
				when "111111111000" => data <= "000000";
				when "111111111001" => data <= "000000";
				when "111111111010" => data <= "000000";
				when "111111111011" => data <= "000000";
				when "111111111100" => data <= "000000";
				when "111111111101" => data <= "000000";
				when "111111111110" => data <= "000000";
				when "111111111111" => data <= "000000";
				when "1000000000000" => data <= "000000";
				when "1000000000001" => data <= "000000";
				when "1000000000010" => data <= "000000";
				when "1000000000011" => data <= "000000";
				when "1000000000100" => data <= "000000";
				when "1000000000101" => data <= "000000";
				when "1000000000110" => data <= "000000";
				when "1000000000111" => data <= "000000";
				when "1000000001000" => data <= "000000";
				when "1000000001001" => data <= "000000";
				when "1000000001010" => data <= "000000";
				when "1000000001011" => data <= "000000";
				when "1000000001100" => data <= "000000";
				when "1000000001101" => data <= "111111";
				when "1000000001110" => data <= "010010";
				when "1000000001111" => data <= "010010";
				when "1000000010000" => data <= "111111";
				when "1000000010001" => data <= "111111";
				when "1000000010010" => data <= "111111";
				when "1000000010011" => data <= "111111";
				when "1000000010100" => data <= "111111";
				when "1000000010101" => data <= "111111";
				when "1000000010110" => data <= "010010";
				when "1000000010111" => data <= "010010";
				when "1000000011000" => data <= "111111";
				when "1000000011001" => data <= "000000";
				when "1000000011010" => data <= "000000";
				when "1000000011011" => data <= "000000";
				when "1000000011100" => data <= "000000";
				when "1000000011101" => data <= "000000";
				when "1000000011110" => data <= "111111";
				when "1000000011111" => data <= "010010";
				when "1000000100000" => data <= "010010";
				when "1000000100001" => data <= "111111";
				when "1000000100010" => data <= "000000";
				when "1000000100011" => data <= "000000";
				when "1000000100100" => data <= "000000";
				when "1000000100101" => data <= "000000";
				when "1000000100110" => data <= "111111";
				when "1000000100111" => data <= "010010";
				when "1000000101000" => data <= "010010";
				when "1000000101001" => data <= "111111";
				when "1000000101010" => data <= "000000";
				when "1000000101011" => data <= "000000";
				when "1000000101100" => data <= "000000";
				when "1000000101101" => data <= "000000";
				when "1000000101110" => data <= "000000";
				when "1000000101111" => data <= "111111";
				when "1000000110000" => data <= "111111";
				when "1000000110001" => data <= "111111";
				when "1000000110010" => data <= "111111";
				when "1000000110011" => data <= "111111";
				when "1000000110100" => data <= "010010";
				when "1000000110101" => data <= "010010";
				when "1000000110110" => data <= "111111";
				when "1000000110111" => data <= "111111";
				when "1000000111000" => data <= "111111";
				when "1000000111001" => data <= "111111";
				when "1000000111010" => data <= "111111";
				when "1000000111011" => data <= "000000";
				when "1000000111100" => data <= "000000";
				when "1000000111101" => data <= "000000";
				when "1000000111110" => data <= "000000";
				when "1000000111111" => data <= "111111";
				when "1000001000000" => data <= "010010";
				when "1000001000001" => data <= "010010";
				when "1000001000010" => data <= "111111";
				when "1000001000011" => data <= "000000";
				when "1000001000100" => data <= "000000";
				when "1000001000101" => data <= "000000";
				when "1000001000110" => data <= "000000";
				when "1000001000111" => data <= "111111";
				when "1000001001000" => data <= "010010";
				when "1000001001001" => data <= "010010";
				when "1000001001010" => data <= "111111";
				when "1000001001011" => data <= "000000";
				when "1000001001100" => data <= "000000";
				when "1000001001101" => data <= "000000";
				when "1000001001110" => data <= "000000";
				when "1000001001111" => data <= "111111";
				when "1000001010000" => data <= "010010";
				when "1000001010001" => data <= "010010";
				when "1000001010010" => data <= "111111";
				when "1000001010011" => data <= "000000";
				when "1000001010100" => data <= "000000";
				when "1000001010101" => data <= "000000";
				when "1000001010110" => data <= "000000";
				when "1000001010111" => data <= "111111";
				when "1000001011000" => data <= "010010";
				when "1000001011001" => data <= "010010";
				when "1000001011010" => data <= "111111";
				when "1000001011011" => data <= "000000";
				when "1000001011100" => data <= "000000";
				when "1000001011101" => data <= "000000";
				when "1000001011110" => data <= "000000";
				when "1000001011111" => data <= "000000";
				when "1000001100000" => data <= "000000";
				when "1000001100001" => data <= "111111";
				when "1000001100010" => data <= "010010";
				when "1000001100011" => data <= "010010";
				when "1000001100100" => data <= "010010";
				when "1000001100101" => data <= "010010";
				when "1000001100110" => data <= "111111";
				when "1000001100111" => data <= "111111";
				when "1000001101000" => data <= "010010";
				when "1000001101001" => data <= "010010";
				when "1000001101010" => data <= "010010";
				when "1000001101011" => data <= "010010";
				when "1000001101100" => data <= "111111";
				when "1000001101101" => data <= "000000";
				when "1000001101110" => data <= "000000";
				when "1000001101111" => data <= "000000";
				when "1000001110000" => data <= "000000";
				when "1000001110001" => data <= "000000";
				when "1000001110010" => data <= "000000";
				when "1000001110011" => data <= "000000";
				when "1000001110100" => data <= "000000";
				when "1000001110101" => data <= "000000";
				when "1000001110110" => data <= "000000";
				when "1000001110111" => data <= "000000";
				when "1000001111000" => data <= "000000";
				when "1000001111001" => data <= "000000";
				when "1000001111010" => data <= "000000";
				when "1000001111011" => data <= "000000";
				when "1000001111100" => data <= "000000";
				when "1000001111101" => data <= "000000";
				when "1000001111110" => data <= "000000";
				when "1000001111111" => data <= "000000";
				when "1000010000000" => data <= "000000";
				when "1000010000001" => data <= "000000";
				when "1000010000010" => data <= "000000";
				when "1000010000011" => data <= "000000";
				when "1000010000100" => data <= "000000";
				when "1000010000101" => data <= "000000";
				when "1000010000110" => data <= "000000";
				when "1000010000111" => data <= "000000";
				when "1000010001000" => data <= "000000";
				when "1000010001001" => data <= "000000";
				when "1000010001010" => data <= "000000";
				when "1000010001011" => data <= "000000";
				when "1000010001100" => data <= "000000";
				when "1000010001101" => data <= "111111";
				when "1000010001110" => data <= "010010";
				when "1000010001111" => data <= "010010";
				when "1000010010000" => data <= "111111";
				when "1000010010001" => data <= "000000";
				when "1000010010010" => data <= "000000";
				when "1000010010011" => data <= "000000";
				when "1000010010100" => data <= "000000";
				when "1000010010101" => data <= "111111";
				when "1000010010110" => data <= "010010";
				when "1000010010111" => data <= "010010";
				when "1000010011000" => data <= "111111";
				when "1000010011001" => data <= "000000";
				when "1000010011010" => data <= "000000";
				when "1000010011011" => data <= "000000";
				when "1000010011100" => data <= "000000";
				when "1000010011101" => data <= "000000";
				when "1000010011110" => data <= "111111";
				when "1000010011111" => data <= "010010";
				when "1000010100000" => data <= "010010";
				when "1000010100001" => data <= "111111";
				when "1000010100010" => data <= "000000";
				when "1000010100011" => data <= "000000";
				when "1000010100100" => data <= "000000";
				when "1000010100101" => data <= "000000";
				when "1000010100110" => data <= "111111";
				when "1000010100111" => data <= "010010";
				when "1000010101000" => data <= "010010";
				when "1000010101001" => data <= "111111";
				when "1000010101010" => data <= "000000";
				when "1000010101011" => data <= "000000";
				when "1000010101100" => data <= "000000";
				when "1000010101101" => data <= "000000";
				when "1000010101110" => data <= "000000";
				when "1000010101111" => data <= "000000";
				when "1000010110000" => data <= "000000";
				when "1000010110001" => data <= "000000";
				when "1000010110010" => data <= "000000";
				when "1000010110011" => data <= "111111";
				when "1000010110100" => data <= "010010";
				when "1000010110101" => data <= "010010";
				when "1000010110110" => data <= "111111";
				when "1000010110111" => data <= "000000";
				when "1000010111000" => data <= "000000";
				when "1000010111001" => data <= "000000";
				when "1000010111010" => data <= "000000";
				when "1000010111011" => data <= "000000";
				when "1000010111100" => data <= "000000";
				when "1000010111101" => data <= "000000";
				when "1000010111110" => data <= "000000";
				when "1000010111111" => data <= "111111";
				when "1000011000000" => data <= "010010";
				when "1000011000001" => data <= "010010";
				when "1000011000010" => data <= "111111";
				when "1000011000011" => data <= "000000";
				when "1000011000100" => data <= "000000";
				when "1000011000101" => data <= "000000";
				when "1000011000110" => data <= "000000";
				when "1000011000111" => data <= "111111";
				when "1000011001000" => data <= "010010";
				when "1000011001001" => data <= "010010";
				when "1000011001010" => data <= "111111";
				when "1000011001011" => data <= "000000";
				when "1000011001100" => data <= "000000";
				when "1000011001101" => data <= "000000";
				when "1000011001110" => data <= "000000";
				when "1000011001111" => data <= "111111";
				when "1000011010000" => data <= "010010";
				when "1000011010001" => data <= "010010";
				when "1000011010010" => data <= "111111";
				when "1000011010011" => data <= "000000";
				when "1000011010100" => data <= "000000";
				when "1000011010101" => data <= "000000";
				when "1000011010110" => data <= "000000";
				when "1000011010111" => data <= "111111";
				when "1000011011000" => data <= "010010";
				when "1000011011001" => data <= "010010";
				when "1000011011010" => data <= "111111";
				when "1000011011011" => data <= "000000";
				when "1000011011100" => data <= "000000";
				when "1000011011101" => data <= "000000";
				when "1000011011110" => data <= "000000";
				when "1000011011111" => data <= "000000";
				when "1000011100000" => data <= "000000";
				when "1000011100001" => data <= "111111";
				when "1000011100010" => data <= "010010";
				when "1000011100011" => data <= "010010";
				when "1000011100100" => data <= "010010";
				when "1000011100101" => data <= "010010";
				when "1000011100110" => data <= "111111";
				when "1000011100111" => data <= "111111";
				when "1000011101000" => data <= "010010";
				when "1000011101001" => data <= "010010";
				when "1000011101010" => data <= "010010";
				when "1000011101011" => data <= "010010";
				when "1000011101100" => data <= "111111";
				when "1000011101101" => data <= "000000";
				when "1000011101110" => data <= "000000";
				when "1000011101111" => data <= "000000";
				when "1000011110000" => data <= "000000";
				when "1000011110001" => data <= "000000";
				when "1000011110010" => data <= "000000";
				when "1000011110011" => data <= "000000";
				when "1000011110100" => data <= "000000";
				when "1000011110101" => data <= "000000";
				when "1000011110110" => data <= "000000";
				when "1000011110111" => data <= "000000";
				when "1000011111000" => data <= "000000";
				when "1000011111001" => data <= "000000";
				when "1000011111010" => data <= "000000";
				when "1000011111011" => data <= "000000";
				when "1000011111100" => data <= "000000";
				when "1000011111101" => data <= "000000";
				when "1000011111110" => data <= "000000";
				when "1000011111111" => data <= "000000";
				when "1000100000000" => data <= "000000";
				when "1000100000001" => data <= "000000";
				when "1000100000010" => data <= "000000";
				when "1000100000011" => data <= "000000";
				when "1000100000100" => data <= "000000";
				when "1000100000101" => data <= "000000";
				when "1000100000110" => data <= "000000";
				when "1000100000111" => data <= "000000";
				when "1000100001000" => data <= "000000";
				when "1000100001001" => data <= "000000";
				when "1000100001010" => data <= "000000";
				when "1000100001011" => data <= "000000";
				when "1000100001100" => data <= "000000";
				when "1000100001101" => data <= "111111";
				when "1000100001110" => data <= "010011";
				when "1000100001111" => data <= "010011";
				when "1000100010000" => data <= "111111";
				when "1000100010001" => data <= "000000";
				when "1000100010010" => data <= "000000";
				when "1000100010011" => data <= "000000";
				when "1000100010100" => data <= "000000";
				when "1000100010101" => data <= "111111";
				when "1000100010110" => data <= "010011";
				when "1000100010111" => data <= "010011";
				when "1000100011000" => data <= "111111";
				when "1000100011001" => data <= "000000";
				when "1000100011010" => data <= "000000";
				when "1000100011011" => data <= "000000";
				when "1000100011100" => data <= "000000";
				when "1000100011101" => data <= "000000";
				when "1000100011110" => data <= "111111";
				when "1000100011111" => data <= "010011";
				when "1000100100000" => data <= "010011";
				when "1000100100001" => data <= "111111";
				when "1000100100010" => data <= "000000";
				when "1000100100011" => data <= "000000";
				when "1000100100100" => data <= "000000";
				when "1000100100101" => data <= "000000";
				when "1000100100110" => data <= "111111";
				when "1000100100111" => data <= "010011";
				when "1000100101000" => data <= "010011";
				when "1000100101001" => data <= "111111";
				when "1000100101010" => data <= "000000";
				when "1000100101011" => data <= "000000";
				when "1000100101100" => data <= "000000";
				when "1000100101101" => data <= "000000";
				when "1000100101110" => data <= "000000";
				when "1000100101111" => data <= "000000";
				when "1000100110000" => data <= "000000";
				when "1000100110001" => data <= "000000";
				when "1000100110010" => data <= "000000";
				when "1000100110011" => data <= "111111";
				when "1000100110100" => data <= "010010";
				when "1000100110101" => data <= "010010";
				when "1000100110110" => data <= "111111";
				when "1000100110111" => data <= "000000";
				when "1000100111000" => data <= "000000";
				when "1000100111001" => data <= "000000";
				when "1000100111010" => data <= "000000";
				when "1000100111011" => data <= "000000";
				when "1000100111100" => data <= "000000";
				when "1000100111101" => data <= "000000";
				when "1000100111110" => data <= "000000";
				when "1000100111111" => data <= "111111";
				when "1000101000000" => data <= "010011";
				when "1000101000001" => data <= "010011";
				when "1000101000010" => data <= "111111";
				when "1000101000011" => data <= "000000";
				when "1000101000100" => data <= "000000";
				when "1000101000101" => data <= "000000";
				when "1000101000110" => data <= "000000";
				when "1000101000111" => data <= "111111";
				when "1000101001000" => data <= "010011";
				when "1000101001001" => data <= "010011";
				when "1000101001010" => data <= "111111";
				when "1000101001011" => data <= "000000";
				when "1000101001100" => data <= "000000";
				when "1000101001101" => data <= "000000";
				when "1000101001110" => data <= "000000";
				when "1000101001111" => data <= "111111";
				when "1000101010000" => data <= "010011";
				when "1000101010001" => data <= "010011";
				when "1000101010010" => data <= "111111";
				when "1000101010011" => data <= "000000";
				when "1000101010100" => data <= "000000";
				when "1000101010101" => data <= "000000";
				when "1000101010110" => data <= "000000";
				when "1000101010111" => data <= "111111";
				when "1000101011000" => data <= "010011";
				when "1000101011001" => data <= "010011";
				when "1000101011010" => data <= "111111";
				when "1000101011011" => data <= "000000";
				when "1000101011100" => data <= "000000";
				when "1000101011101" => data <= "000000";
				when "1000101011110" => data <= "000000";
				when "1000101011111" => data <= "000000";
				when "1000101100000" => data <= "000000";
				when "1000101100001" => data <= "111111";
				when "1000101100010" => data <= "010010";
				when "1000101100011" => data <= "010010";
				when "1000101100100" => data <= "111111";
				when "1000101100101" => data <= "111111";
				when "1000101100110" => data <= "010010";
				when "1000101100111" => data <= "010010";
				when "1000101101000" => data <= "111111";
				when "1000101101001" => data <= "111111";
				when "1000101101010" => data <= "010010";
				when "1000101101011" => data <= "010010";
				when "1000101101100" => data <= "111111";
				when "1000101101101" => data <= "000000";
				when "1000101101110" => data <= "000000";
				when "1000101101111" => data <= "000000";
				when "1000101110000" => data <= "000000";
				when "1000101110001" => data <= "000000";
				when "1000101110010" => data <= "000000";
				when "1000101110011" => data <= "000000";
				when "1000101110100" => data <= "000000";
				when "1000101110101" => data <= "000000";
				when "1000101110110" => data <= "000000";
				when "1000101110111" => data <= "000000";
				when "1000101111000" => data <= "000000";
				when "1000101111001" => data <= "000000";
				when "1000101111010" => data <= "000000";
				when "1000101111011" => data <= "000000";
				when "1000101111100" => data <= "000000";
				when "1000101111101" => data <= "000000";
				when "1000101111110" => data <= "000000";
				when "1000101111111" => data <= "000000";
				when "1000110000000" => data <= "000000";
				when "1000110000001" => data <= "000000";
				when "1000110000010" => data <= "000000";
				when "1000110000011" => data <= "000000";
				when "1000110000100" => data <= "000000";
				when "1000110000101" => data <= "000000";
				when "1000110000110" => data <= "000000";
				when "1000110000111" => data <= "000000";
				when "1000110001000" => data <= "000000";
				when "1000110001001" => data <= "000000";
				when "1000110001010" => data <= "000000";
				when "1000110001011" => data <= "000000";
				when "1000110001100" => data <= "000000";
				when "1000110001101" => data <= "111111";
				when "1000110001110" => data <= "010011";
				when "1000110001111" => data <= "010011";
				when "1000110010000" => data <= "111111";
				when "1000110010001" => data <= "000000";
				when "1000110010010" => data <= "000000";
				when "1000110010011" => data <= "000000";
				when "1000110010100" => data <= "000000";
				when "1000110010101" => data <= "111111";
				when "1000110010110" => data <= "010011";
				when "1000110010111" => data <= "010011";
				when "1000110011000" => data <= "111111";
				when "1000110011001" => data <= "000000";
				when "1000110011010" => data <= "000000";
				when "1000110011011" => data <= "000000";
				when "1000110011100" => data <= "000000";
				when "1000110011101" => data <= "000000";
				when "1000110011110" => data <= "111111";
				when "1000110011111" => data <= "010011";
				when "1000110100000" => data <= "010011";
				when "1000110100001" => data <= "111111";
				when "1000110100010" => data <= "111111";
				when "1000110100011" => data <= "000000";
				when "1000110100100" => data <= "000000";
				when "1000110100101" => data <= "111111";
				when "1000110100110" => data <= "111111";
				when "1000110100111" => data <= "010011";
				when "1000110101000" => data <= "010011";
				when "1000110101001" => data <= "111111";
				when "1000110101010" => data <= "000000";
				when "1000110101011" => data <= "000000";
				when "1000110101100" => data <= "000000";
				when "1000110101101" => data <= "000000";
				when "1000110101110" => data <= "000000";
				when "1000110101111" => data <= "000000";
				when "1000110110000" => data <= "000000";
				when "1000110110001" => data <= "000000";
				when "1000110110010" => data <= "000000";
				when "1000110110011" => data <= "111111";
				when "1000110110100" => data <= "010011";
				when "1000110110101" => data <= "010011";
				when "1000110110110" => data <= "111111";
				when "1000110110111" => data <= "000000";
				when "1000110111000" => data <= "000000";
				when "1000110111001" => data <= "000000";
				when "1000110111010" => data <= "000000";
				when "1000110111011" => data <= "000000";
				when "1000110111100" => data <= "000000";
				when "1000110111101" => data <= "000000";
				when "1000110111110" => data <= "000000";
				when "1000110111111" => data <= "111111";
				when "1000111000000" => data <= "010011";
				when "1000111000001" => data <= "010011";
				when "1000111000010" => data <= "111111";
				when "1000111000011" => data <= "000000";
				when "1000111000100" => data <= "000000";
				when "1000111000101" => data <= "000000";
				when "1000111000110" => data <= "000000";
				when "1000111000111" => data <= "111111";
				when "1000111001000" => data <= "010011";
				when "1000111001001" => data <= "010011";
				when "1000111001010" => data <= "111111";
				when "1000111001011" => data <= "000000";
				when "1000111001100" => data <= "000000";
				when "1000111001101" => data <= "000000";
				when "1000111001110" => data <= "000000";
				when "1000111001111" => data <= "111111";
				when "1000111010000" => data <= "010011";
				when "1000111010001" => data <= "010011";
				when "1000111010010" => data <= "111111";
				when "1000111010011" => data <= "111111";
				when "1000111010100" => data <= "000000";
				when "1000111010101" => data <= "000000";
				when "1000111010110" => data <= "111111";
				when "1000111010111" => data <= "111111";
				when "1000111011000" => data <= "010011";
				when "1000111011001" => data <= "010011";
				when "1000111011010" => data <= "111111";
				when "1000111011011" => data <= "000000";
				when "1000111011100" => data <= "000000";
				when "1000111011101" => data <= "000000";
				when "1000111011110" => data <= "000000";
				when "1000111011111" => data <= "000000";
				when "1000111100000" => data <= "000000";
				when "1000111100001" => data <= "111111";
				when "1000111100010" => data <= "010010";
				when "1000111100011" => data <= "010010";
				when "1000111100100" => data <= "111111";
				when "1000111100101" => data <= "111111";
				when "1000111100110" => data <= "010010";
				when "1000111100111" => data <= "010010";
				when "1000111101000" => data <= "111111";
				when "1000111101001" => data <= "111111";
				when "1000111101010" => data <= "010010";
				when "1000111101011" => data <= "010010";
				when "1000111101100" => data <= "111111";
				when "1000111101101" => data <= "000000";
				when "1000111101110" => data <= "000000";
				when "1000111101111" => data <= "000000";
				when "1000111110000" => data <= "000000";
				when "1000111110001" => data <= "000000";
				when "1000111110010" => data <= "000000";
				when "1000111110011" => data <= "000000";
				when "1000111110100" => data <= "000000";
				when "1000111110101" => data <= "000000";
				when "1000111110110" => data <= "000000";
				when "1000111110111" => data <= "000000";
				when "1000111111000" => data <= "000000";
				when "1000111111001" => data <= "000000";
				when "1000111111010" => data <= "000000";
				when "1000111111011" => data <= "000000";
				when "1000111111100" => data <= "000000";
				when "1000111111101" => data <= "000000";
				when "1000111111110" => data <= "000000";
				when "1000111111111" => data <= "000000";
				when "1001000000000" => data <= "000000";
				when "1001000000001" => data <= "000000";
				when "1001000000010" => data <= "000000";
				when "1001000000011" => data <= "000000";
				when "1001000000100" => data <= "000000";
				when "1001000000101" => data <= "000000";
				when "1001000000110" => data <= "000000";
				when "1001000000111" => data <= "000000";
				when "1001000001000" => data <= "000000";
				when "1001000001001" => data <= "000000";
				when "1001000001010" => data <= "000000";
				when "1001000001011" => data <= "000000";
				when "1001000001100" => data <= "000000";
				when "1001000001101" => data <= "111111";
				when "1001000001110" => data <= "010011";
				when "1001000001111" => data <= "010011";
				when "1001000010000" => data <= "111111";
				when "1001000010001" => data <= "000000";
				when "1001000010010" => data <= "000000";
				when "1001000010011" => data <= "000000";
				when "1001000010100" => data <= "000000";
				when "1001000010101" => data <= "111111";
				when "1001000010110" => data <= "010011";
				when "1001000010111" => data <= "010011";
				when "1001000011000" => data <= "111111";
				when "1001000011001" => data <= "000000";
				when "1001000011010" => data <= "000000";
				when "1001000011011" => data <= "000000";
				when "1001000011100" => data <= "000000";
				when "1001000011101" => data <= "000000";
				when "1001000011110" => data <= "000000";
				when "1001000011111" => data <= "111111";
				when "1001000100000" => data <= "111111";
				when "1001000100001" => data <= "010011";
				when "1001000100010" => data <= "010011";
				when "1001000100011" => data <= "111111";
				when "1001000100100" => data <= "111111";
				when "1001000100101" => data <= "010011";
				when "1001000100110" => data <= "010011";
				when "1001000100111" => data <= "111111";
				when "1001000101000" => data <= "111111";
				when "1001000101001" => data <= "000000";
				when "1001000101010" => data <= "000000";
				when "1001000101011" => data <= "000000";
				when "1001000101100" => data <= "000000";
				when "1001000101101" => data <= "000000";
				when "1001000101110" => data <= "000000";
				when "1001000101111" => data <= "000000";
				when "1001000110000" => data <= "000000";
				when "1001000110001" => data <= "000000";
				when "1001000110010" => data <= "000000";
				when "1001000110011" => data <= "111111";
				when "1001000110100" => data <= "010011";
				when "1001000110101" => data <= "010011";
				when "1001000110110" => data <= "111111";
				when "1001000110111" => data <= "000000";
				when "1001000111000" => data <= "000000";
				when "1001000111001" => data <= "000000";
				when "1001000111010" => data <= "000000";
				when "1001000111011" => data <= "000000";
				when "1001000111100" => data <= "000000";
				when "1001000111101" => data <= "000000";
				when "1001000111110" => data <= "000000";
				when "1001000111111" => data <= "111111";
				when "1001001000000" => data <= "010011";
				when "1001001000001" => data <= "010011";
				when "1001001000010" => data <= "111111";
				when "1001001000011" => data <= "111111";
				when "1001001000100" => data <= "111111";
				when "1001001000101" => data <= "111111";
				when "1001001000110" => data <= "111111";
				when "1001001000111" => data <= "111111";
				when "1001001001000" => data <= "010011";
				when "1001001001001" => data <= "010011";
				when "1001001001010" => data <= "111111";
				when "1001001001011" => data <= "000000";
				when "1001001001100" => data <= "000000";
				when "1001001001101" => data <= "000000";
				when "1001001001110" => data <= "000000";
				when "1001001001111" => data <= "000000";
				when "1001001010000" => data <= "111111";
				when "1001001010001" => data <= "111111";
				when "1001001010010" => data <= "010011";
				when "1001001010011" => data <= "010011";
				when "1001001010100" => data <= "111111";
				when "1001001010101" => data <= "111111";
				when "1001001010110" => data <= "010011";
				when "1001001010111" => data <= "010011";
				when "1001001011000" => data <= "111111";
				when "1001001011001" => data <= "111111";
				when "1001001011010" => data <= "000000";
				when "1001001011011" => data <= "000000";
				when "1001001011100" => data <= "000000";
				when "1001001011101" => data <= "000000";
				when "1001001011110" => data <= "000000";
				when "1001001011111" => data <= "000000";
				when "1001001100000" => data <= "000000";
				when "1001001100001" => data <= "111111";
				when "1001001100010" => data <= "010011";
				when "1001001100011" => data <= "010011";
				when "1001001100100" => data <= "111111";
				when "1001001100101" => data <= "000000";
				when "1001001100110" => data <= "111111";
				when "1001001100111" => data <= "111111";
				when "1001001101000" => data <= "000000";
				when "1001001101001" => data <= "111111";
				when "1001001101010" => data <= "010011";
				when "1001001101011" => data <= "010011";
				when "1001001101100" => data <= "111111";
				when "1001001101101" => data <= "000000";
				when "1001001101110" => data <= "000000";
				when "1001001101111" => data <= "000000";
				when "1001001110000" => data <= "000000";
				when "1001001110001" => data <= "000000";
				when "1001001110010" => data <= "000000";
				when "1001001110011" => data <= "000000";
				when "1001001110100" => data <= "000000";
				when "1001001110101" => data <= "000000";
				when "1001001110110" => data <= "000000";
				when "1001001110111" => data <= "000000";
				when "1001001111000" => data <= "000000";
				when "1001001111001" => data <= "000000";
				when "1001001111010" => data <= "000000";
				when "1001001111011" => data <= "000000";
				when "1001001111100" => data <= "000000";
				when "1001001111101" => data <= "000000";
				when "1001001111110" => data <= "000000";
				when "1001001111111" => data <= "000000";
				when "1001010000000" => data <= "000000";
				when "1001010000001" => data <= "000000";
				when "1001010000010" => data <= "000000";
				when "1001010000011" => data <= "000000";
				when "1001010000100" => data <= "000000";
				when "1001010000101" => data <= "000000";
				when "1001010000110" => data <= "000000";
				when "1001010000111" => data <= "000000";
				when "1001010001000" => data <= "000000";
				when "1001010001001" => data <= "000000";
				when "1001010001010" => data <= "000000";
				when "1001010001011" => data <= "000000";
				when "1001010001100" => data <= "000000";
				when "1001010001101" => data <= "111111";
				when "1001010001110" => data <= "010011";
				when "1001010001111" => data <= "010011";
				when "1001010010000" => data <= "111111";
				when "1001010010001" => data <= "111111";
				when "1001010010010" => data <= "111111";
				when "1001010010011" => data <= "111111";
				when "1001010010100" => data <= "111111";
				when "1001010010101" => data <= "111111";
				when "1001010010110" => data <= "010011";
				when "1001010010111" => data <= "010011";
				when "1001010011000" => data <= "111111";
				when "1001010011001" => data <= "000000";
				when "1001010011010" => data <= "000000";
				when "1001010011011" => data <= "000000";
				when "1001010011100" => data <= "000000";
				when "1001010011101" => data <= "000000";
				when "1001010011110" => data <= "000000";
				when "1001010011111" => data <= "000000";
				when "1001010100000" => data <= "111111";
				when "1001010100001" => data <= "010011";
				when "1001010100010" => data <= "010011";
				when "1001010100011" => data <= "111111";
				when "1001010100100" => data <= "111111";
				when "1001010100101" => data <= "010011";
				when "1001010100110" => data <= "010011";
				when "1001010100111" => data <= "111111";
				when "1001010101000" => data <= "000000";
				when "1001010101001" => data <= "000000";
				when "1001010101010" => data <= "000000";
				when "1001010101011" => data <= "000000";
				when "1001010101100" => data <= "000000";
				when "1001010101101" => data <= "000000";
				when "1001010101110" => data <= "000000";
				when "1001010101111" => data <= "000000";
				when "1001010110000" => data <= "000000";
				when "1001010110001" => data <= "000000";
				when "1001010110010" => data <= "000000";
				when "1001010110011" => data <= "111111";
				when "1001010110100" => data <= "010011";
				when "1001010110101" => data <= "010011";
				when "1001010110110" => data <= "111111";
				when "1001010110111" => data <= "000000";
				when "1001010111000" => data <= "000000";
				when "1001010111001" => data <= "000000";
				when "1001010111010" => data <= "000000";
				when "1001010111011" => data <= "000000";
				when "1001010111100" => data <= "000000";
				when "1001010111101" => data <= "000000";
				when "1001010111110" => data <= "000000";
				when "1001010111111" => data <= "111111";
				when "1001011000000" => data <= "010011";
				when "1001011000001" => data <= "010011";
				when "1001011000010" => data <= "010011";
				when "1001011000011" => data <= "010011";
				when "1001011000100" => data <= "010011";
				when "1001011000101" => data <= "010011";
				when "1001011000110" => data <= "010011";
				when "1001011000111" => data <= "010011";
				when "1001011001000" => data <= "010011";
				when "1001011001001" => data <= "010011";
				when "1001011001010" => data <= "111111";
				when "1001011001011" => data <= "000000";
				when "1001011001100" => data <= "000000";
				when "1001011001101" => data <= "000000";
				when "1001011001110" => data <= "000000";
				when "1001011001111" => data <= "000000";
				when "1001011010000" => data <= "000000";
				when "1001011010001" => data <= "111111";
				when "1001011010010" => data <= "010011";
				when "1001011010011" => data <= "010011";
				when "1001011010100" => data <= "111111";
				when "1001011010101" => data <= "111111";
				when "1001011010110" => data <= "010011";
				when "1001011010111" => data <= "010011";
				when "1001011011000" => data <= "111111";
				when "1001011011001" => data <= "000000";
				when "1001011011010" => data <= "000000";
				when "1001011011011" => data <= "000000";
				when "1001011011100" => data <= "000000";
				when "1001011011101" => data <= "000000";
				when "1001011011110" => data <= "000000";
				when "1001011011111" => data <= "000000";
				when "1001011100000" => data <= "000000";
				when "1001011100001" => data <= "111111";
				when "1001011100010" => data <= "010011";
				when "1001011100011" => data <= "010011";
				when "1001011100100" => data <= "111111";
				when "1001011100101" => data <= "000000";
				when "1001011100110" => data <= "000000";
				when "1001011100111" => data <= "000000";
				when "1001011101000" => data <= "000000";
				when "1001011101001" => data <= "111111";
				when "1001011101010" => data <= "010011";
				when "1001011101011" => data <= "010011";
				when "1001011101100" => data <= "111111";
				when "1001011101101" => data <= "000000";
				when "1001011101110" => data <= "000000";
				when "1001011101111" => data <= "000000";
				when "1001011110000" => data <= "000000";
				when "1001011110001" => data <= "000000";
				when "1001011110010" => data <= "000000";
				when "1001011110011" => data <= "000000";
				when "1001011110100" => data <= "000000";
				when "1001011110101" => data <= "000000";
				when "1001011110110" => data <= "000000";
				when "1001011110111" => data <= "000000";
				when "1001011111000" => data <= "000000";
				when "1001011111001" => data <= "000000";
				when "1001011111010" => data <= "000000";
				when "1001011111011" => data <= "000000";
				when "1001011111100" => data <= "000000";
				when "1001011111101" => data <= "000000";
				when "1001011111110" => data <= "000000";
				when "1001011111111" => data <= "000000";
				when "1001100000000" => data <= "000000";
				when "1001100000001" => data <= "000000";
				when "1001100000010" => data <= "000000";
				when "1001100000011" => data <= "000000";
				when "1001100000100" => data <= "000000";
				when "1001100000101" => data <= "000000";
				when "1001100000110" => data <= "000000";
				when "1001100000111" => data <= "000000";
				when "1001100001000" => data <= "000000";
				when "1001100001001" => data <= "000000";
				when "1001100001010" => data <= "000000";
				when "1001100001011" => data <= "000000";
				when "1001100001100" => data <= "000000";
				when "1001100001101" => data <= "111111";
				when "1001100001110" => data <= "010011";
				when "1001100001111" => data <= "010011";
				when "1001100010000" => data <= "010011";
				when "1001100010001" => data <= "010011";
				when "1001100010010" => data <= "010011";
				when "1001100010011" => data <= "010011";
				when "1001100010100" => data <= "010011";
				when "1001100010101" => data <= "010011";
				when "1001100010110" => data <= "111111";
				when "1001100010111" => data <= "111111";
				when "1001100011000" => data <= "000000";
				when "1001100011001" => data <= "000000";
				when "1001100011010" => data <= "000000";
				when "1001100011011" => data <= "000000";
				when "1001100011100" => data <= "000000";
				when "1001100011101" => data <= "000000";
				when "1001100011110" => data <= "000000";
				when "1001100011111" => data <= "000000";
				when "1001100100000" => data <= "000000";
				when "1001100100001" => data <= "111111";
				when "1001100100010" => data <= "111111";
				when "1001100100011" => data <= "010011";
				when "1001100100100" => data <= "010011";
				when "1001100100101" => data <= "111111";
				when "1001100100110" => data <= "111111";
				when "1001100100111" => data <= "000000";
				when "1001100101000" => data <= "000000";
				when "1001100101001" => data <= "000000";
				when "1001100101010" => data <= "000000";
				when "1001100101011" => data <= "000000";
				when "1001100101100" => data <= "000000";
				when "1001100101101" => data <= "000000";
				when "1001100101110" => data <= "000000";
				when "1001100101111" => data <= "000000";
				when "1001100110000" => data <= "000000";
				when "1001100110001" => data <= "000000";
				when "1001100110010" => data <= "000000";
				when "1001100110011" => data <= "111111";
				when "1001100110100" => data <= "010011";
				when "1001100110101" => data <= "010011";
				when "1001100110110" => data <= "111111";
				when "1001100110111" => data <= "000000";
				when "1001100111000" => data <= "000000";
				when "1001100111001" => data <= "000000";
				when "1001100111010" => data <= "000000";
				when "1001100111011" => data <= "000000";
				when "1001100111100" => data <= "000000";
				when "1001100111101" => data <= "000000";
				when "1001100111110" => data <= "000000";
				when "1001100111111" => data <= "111111";
				when "1001101000000" => data <= "010011";
				when "1001101000001" => data <= "010011";
				when "1001101000010" => data <= "010011";
				when "1001101000011" => data <= "010011";
				when "1001101000100" => data <= "010011";
				when "1001101000101" => data <= "010011";
				when "1001101000110" => data <= "010011";
				when "1001101000111" => data <= "010011";
				when "1001101001000" => data <= "010011";
				when "1001101001001" => data <= "010011";
				when "1001101001010" => data <= "111111";
				when "1001101001011" => data <= "000000";
				when "1001101001100" => data <= "000000";
				when "1001101001101" => data <= "000000";
				when "1001101001110" => data <= "000000";
				when "1001101001111" => data <= "000000";
				when "1001101010000" => data <= "000000";
				when "1001101010001" => data <= "000000";
				when "1001101010010" => data <= "111111";
				when "1001101010011" => data <= "111111";
				when "1001101010100" => data <= "010011";
				when "1001101010101" => data <= "010011";
				when "1001101010110" => data <= "111111";
				when "1001101010111" => data <= "111111";
				when "1001101011000" => data <= "000000";
				when "1001101011001" => data <= "000000";
				when "1001101011010" => data <= "000000";
				when "1001101011011" => data <= "000000";
				when "1001101011100" => data <= "000000";
				when "1001101011101" => data <= "000000";
				when "1001101011110" => data <= "000000";
				when "1001101011111" => data <= "000000";
				when "1001101100000" => data <= "000000";
				when "1001101100001" => data <= "111111";
				when "1001101100010" => data <= "010011";
				when "1001101100011" => data <= "010011";
				when "1001101100100" => data <= "111111";
				when "1001101100101" => data <= "000000";
				when "1001101100110" => data <= "000000";
				when "1001101100111" => data <= "000000";
				when "1001101101000" => data <= "000000";
				when "1001101101001" => data <= "111111";
				when "1001101101010" => data <= "010011";
				when "1001101101011" => data <= "010011";
				when "1001101101100" => data <= "111111";
				when "1001101101101" => data <= "000000";
				when "1001101101110" => data <= "000000";
				when "1001101101111" => data <= "000000";
				when "1001101110000" => data <= "000000";
				when "1001101110001" => data <= "000000";
				when "1001101110010" => data <= "000000";
				when "1001101110011" => data <= "000000";
				when "1001101110100" => data <= "000000";
				when "1001101110101" => data <= "000000";
				when "1001101110110" => data <= "000000";
				when "1001101110111" => data <= "000000";
				when "1001101111000" => data <= "000000";
				when "1001101111001" => data <= "000000";
				when "1001101111010" => data <= "000000";
				when "1001101111011" => data <= "000000";
				when "1001101111100" => data <= "000000";
				when "1001101111101" => data <= "000000";
				when "1001101111110" => data <= "000000";
				when "1001101111111" => data <= "000000";
				when "1001110000000" => data <= "000000";
				when "1001110000001" => data <= "000000";
				when "1001110000010" => data <= "000000";
				when "1001110000011" => data <= "000000";
				when "1001110000100" => data <= "000000";
				when "1001110000101" => data <= "000000";
				when "1001110000110" => data <= "000000";
				when "1001110000111" => data <= "000000";
				when "1001110001000" => data <= "000000";
				when "1001110001001" => data <= "000000";
				when "1001110001010" => data <= "000000";
				when "1001110001011" => data <= "000000";
				when "1001110001100" => data <= "000000";
				when "1001110001101" => data <= "111111";
				when "1001110001110" => data <= "010011";
				when "1001110001111" => data <= "010011";
				when "1001110010000" => data <= "010011";
				when "1001110010001" => data <= "010011";
				when "1001110010010" => data <= "010011";
				when "1001110010011" => data <= "010011";
				when "1001110010100" => data <= "010011";
				when "1001110010101" => data <= "010011";
				when "1001110010110" => data <= "111111";
				when "1001110010111" => data <= "000000";
				when "1001110011000" => data <= "000000";
				when "1001110011001" => data <= "000000";
				when "1001110011010" => data <= "000000";
				when "1001110011011" => data <= "000000";
				when "1001110011100" => data <= "000000";
				when "1001110011101" => data <= "000000";
				when "1001110011110" => data <= "000000";
				when "1001110011111" => data <= "000000";
				when "1001110100000" => data <= "000000";
				when "1001110100001" => data <= "000000";
				when "1001110100010" => data <= "111111";
				when "1001110100011" => data <= "010011";
				when "1001110100100" => data <= "010011";
				when "1001110100101" => data <= "111111";
				when "1001110100110" => data <= "000000";
				when "1001110100111" => data <= "000000";
				when "1001110101000" => data <= "000000";
				when "1001110101001" => data <= "000000";
				when "1001110101010" => data <= "000000";
				when "1001110101011" => data <= "000000";
				when "1001110101100" => data <= "000000";
				when "1001110101101" => data <= "000000";
				when "1001110101110" => data <= "000000";
				when "1001110101111" => data <= "000000";
				when "1001110110000" => data <= "000000";
				when "1001110110001" => data <= "000000";
				when "1001110110010" => data <= "000000";
				when "1001110110011" => data <= "111111";
				when "1001110110100" => data <= "010011";
				when "1001110110101" => data <= "010011";
				when "1001110110110" => data <= "111111";
				when "1001110110111" => data <= "000000";
				when "1001110111000" => data <= "000000";
				when "1001110111001" => data <= "000000";
				when "1001110111010" => data <= "000000";
				when "1001110111011" => data <= "000000";
				when "1001110111100" => data <= "000000";
				when "1001110111101" => data <= "000000";
				when "1001110111110" => data <= "000000";
				when "1001110111111" => data <= "111111";
				when "1001111000000" => data <= "010011";
				when "1001111000001" => data <= "010011";
				when "1001111000010" => data <= "111111";
				when "1001111000011" => data <= "111111";
				when "1001111000100" => data <= "111111";
				when "1001111000101" => data <= "111111";
				when "1001111000110" => data <= "111111";
				when "1001111000111" => data <= "111111";
				when "1001111001000" => data <= "010011";
				when "1001111001001" => data <= "010011";
				when "1001111001010" => data <= "111111";
				when "1001111001011" => data <= "000000";
				when "1001111001100" => data <= "000000";
				when "1001111001101" => data <= "000000";
				when "1001111001110" => data <= "000000";
				when "1001111001111" => data <= "000000";
				when "1001111010000" => data <= "000000";
				when "1001111010001" => data <= "000000";
				when "1001111010010" => data <= "000000";
				when "1001111010011" => data <= "111111";
				when "1001111010100" => data <= "010011";
				when "1001111010101" => data <= "010011";
				when "1001111010110" => data <= "111111";
				when "1001111010111" => data <= "000000";
				when "1001111011000" => data <= "000000";
				when "1001111011001" => data <= "000000";
				when "1001111011010" => data <= "000000";
				when "1001111011011" => data <= "000000";
				when "1001111011100" => data <= "000000";
				when "1001111011101" => data <= "000000";
				when "1001111011110" => data <= "000000";
				when "1001111011111" => data <= "000000";
				when "1001111100000" => data <= "000000";
				when "1001111100001" => data <= "111111";
				when "1001111100010" => data <= "100011";
				when "1001111100011" => data <= "100011";
				when "1001111100100" => data <= "111111";
				when "1001111100101" => data <= "000000";
				when "1001111100110" => data <= "000000";
				when "1001111100111" => data <= "000000";
				when "1001111101000" => data <= "000000";
				when "1001111101001" => data <= "111111";
				when "1001111101010" => data <= "100011";
				when "1001111101011" => data <= "100011";
				when "1001111101100" => data <= "111111";
				when "1001111101101" => data <= "000000";
				when "1001111101110" => data <= "000000";
				when "1001111101111" => data <= "000000";
				when "1001111110000" => data <= "000000";
				when "1001111110001" => data <= "000000";
				when "1001111110010" => data <= "000000";
				when "1001111110011" => data <= "000000";
				when "1001111110100" => data <= "000000";
				when "1001111110101" => data <= "000000";
				when "1001111110110" => data <= "000000";
				when "1001111110111" => data <= "000000";
				when "1001111111000" => data <= "000000";
				when "1001111111001" => data <= "000000";
				when "1001111111010" => data <= "000000";
				when "1001111111011" => data <= "000000";
				when "1001111111100" => data <= "000000";
				when "1001111111101" => data <= "000000";
				when "1001111111110" => data <= "000000";
				when "1001111111111" => data <= "000000";
				when "1010000000000" => data <= "000000";
				when "1010000000001" => data <= "000000";
				when "1010000000010" => data <= "000000";
				when "1010000000011" => data <= "000000";
				when "1010000000100" => data <= "000000";
				when "1010000000101" => data <= "000000";
				when "1010000000110" => data <= "000000";
				when "1010000000111" => data <= "000000";
				when "1010000001000" => data <= "000000";
				when "1010000001001" => data <= "000000";
				when "1010000001010" => data <= "000000";
				when "1010000001011" => data <= "000000";
				when "1010000001100" => data <= "000000";
				when "1010000001101" => data <= "111111";
				when "1010000001110" => data <= "100011";
				when "1010000001111" => data <= "100011";
				when "1010000010000" => data <= "111111";
				when "1010000010001" => data <= "111111";
				when "1010000010010" => data <= "111111";
				when "1010000010011" => data <= "111111";
				when "1010000010100" => data <= "111111";
				when "1010000010101" => data <= "111111";
				when "1010000010110" => data <= "100011";
				when "1010000010111" => data <= "111111";
				when "1010000011000" => data <= "000000";
				when "1010000011001" => data <= "000000";
				when "1010000011010" => data <= "000000";
				when "1010000011011" => data <= "000000";
				when "1010000011100" => data <= "000000";
				when "1010000011101" => data <= "000000";
				when "1010000011110" => data <= "000000";
				when "1010000011111" => data <= "000000";
				when "1010000100000" => data <= "000000";
				when "1010000100001" => data <= "000000";
				when "1010000100010" => data <= "111111";
				when "1010000100011" => data <= "100011";
				when "1010000100100" => data <= "100011";
				when "1010000100101" => data <= "111111";
				when "1010000100110" => data <= "000000";
				when "1010000100111" => data <= "000000";
				when "1010000101000" => data <= "000000";
				when "1010000101001" => data <= "000000";
				when "1010000101010" => data <= "000000";
				when "1010000101011" => data <= "000000";
				when "1010000101100" => data <= "000000";
				when "1010000101101" => data <= "000000";
				when "1010000101110" => data <= "000000";
				when "1010000101111" => data <= "000000";
				when "1010000110000" => data <= "000000";
				when "1010000110001" => data <= "000000";
				when "1010000110010" => data <= "000000";
				when "1010000110011" => data <= "111111";
				when "1010000110100" => data <= "100011";
				when "1010000110101" => data <= "100011";
				when "1010000110110" => data <= "111111";
				when "1010000110111" => data <= "000000";
				when "1010000111000" => data <= "000000";
				when "1010000111001" => data <= "000000";
				when "1010000111010" => data <= "000000";
				when "1010000111011" => data <= "000000";
				when "1010000111100" => data <= "000000";
				when "1010000111101" => data <= "000000";
				when "1010000111110" => data <= "000000";
				when "1010000111111" => data <= "111111";
				when "1010001000000" => data <= "100011";
				when "1010001000001" => data <= "100011";
				when "1010001000010" => data <= "111111";
				when "1010001000011" => data <= "000000";
				when "1010001000100" => data <= "000000";
				when "1010001000101" => data <= "000000";
				when "1010001000110" => data <= "000000";
				when "1010001000111" => data <= "111111";
				when "1010001001000" => data <= "100011";
				when "1010001001001" => data <= "100011";
				when "1010001001010" => data <= "111111";
				when "1010001001011" => data <= "000000";
				when "1010001001100" => data <= "000000";
				when "1010001001101" => data <= "000000";
				when "1010001001110" => data <= "000000";
				when "1010001001111" => data <= "000000";
				when "1010001010000" => data <= "000000";
				when "1010001010001" => data <= "000000";
				when "1010001010010" => data <= "000000";
				when "1010001010011" => data <= "111111";
				when "1010001010100" => data <= "100011";
				when "1010001010101" => data <= "100011";
				when "1010001010110" => data <= "111111";
				when "1010001010111" => data <= "000000";
				when "1010001011000" => data <= "000000";
				when "1010001011001" => data <= "000000";
				when "1010001011010" => data <= "000000";
				when "1010001011011" => data <= "000000";
				when "1010001011100" => data <= "000000";
				when "1010001011101" => data <= "000000";
				when "1010001011110" => data <= "000000";
				when "1010001011111" => data <= "000000";
				when "1010001100000" => data <= "000000";
				when "1010001100001" => data <= "111111";
				when "1010001100010" => data <= "100011";
				when "1010001100011" => data <= "100011";
				when "1010001100100" => data <= "111111";
				when "1010001100101" => data <= "000000";
				when "1010001100110" => data <= "000000";
				when "1010001100111" => data <= "000000";
				when "1010001101000" => data <= "000000";
				when "1010001101001" => data <= "111111";
				when "1010001101010" => data <= "100011";
				when "1010001101011" => data <= "100011";
				when "1010001101100" => data <= "111111";
				when "1010001101101" => data <= "000000";
				when "1010001101110" => data <= "000000";
				when "1010001101111" => data <= "000000";
				when "1010001110000" => data <= "000000";
				when "1010001110001" => data <= "000000";
				when "1010001110010" => data <= "000000";
				when "1010001110011" => data <= "000000";
				when "1010001110100" => data <= "000000";
				when "1010001110101" => data <= "000000";
				when "1010001110110" => data <= "000000";
				when "1010001110111" => data <= "000000";
				when "1010001111000" => data <= "000000";
				when "1010001111001" => data <= "000000";
				when "1010001111010" => data <= "000000";
				when "1010001111011" => data <= "000000";
				when "1010001111100" => data <= "000000";
				when "1010001111101" => data <= "000000";
				when "1010001111110" => data <= "000000";
				when "1010001111111" => data <= "000000";
				when "1010010000000" => data <= "000000";
				when "1010010000001" => data <= "000000";
				when "1010010000010" => data <= "000000";
				when "1010010000011" => data <= "000000";
				when "1010010000100" => data <= "000000";
				when "1010010000101" => data <= "000000";
				when "1010010000110" => data <= "000000";
				when "1010010000111" => data <= "000000";
				when "1010010001000" => data <= "000000";
				when "1010010001001" => data <= "000000";
				when "1010010001010" => data <= "000000";
				when "1010010001011" => data <= "000000";
				when "1010010001100" => data <= "000000";
				when "1010010001101" => data <= "111111";
				when "1010010001110" => data <= "100011";
				when "1010010001111" => data <= "100011";
				when "1010010010000" => data <= "111111";
				when "1010010010001" => data <= "000000";
				when "1010010010010" => data <= "000000";
				when "1010010010011" => data <= "000000";
				when "1010010010100" => data <= "000000";
				when "1010010010101" => data <= "111111";
				when "1010010010110" => data <= "100011";
				when "1010010010111" => data <= "100011";
				when "1010010011000" => data <= "111111";
				when "1010010011001" => data <= "000000";
				when "1010010011010" => data <= "000000";
				when "1010010011011" => data <= "000000";
				when "1010010011100" => data <= "000000";
				when "1010010011101" => data <= "000000";
				when "1010010011110" => data <= "000000";
				when "1010010011111" => data <= "000000";
				when "1010010100000" => data <= "000000";
				when "1010010100001" => data <= "000000";
				when "1010010100010" => data <= "111111";
				when "1010010100011" => data <= "100011";
				when "1010010100100" => data <= "100011";
				when "1010010100101" => data <= "111111";
				when "1010010100110" => data <= "000000";
				when "1010010100111" => data <= "000000";
				when "1010010101000" => data <= "000000";
				when "1010010101001" => data <= "000000";
				when "1010010101010" => data <= "000000";
				when "1010010101011" => data <= "000000";
				when "1010010101100" => data <= "000000";
				when "1010010101101" => data <= "000000";
				when "1010010101110" => data <= "000000";
				when "1010010101111" => data <= "000000";
				when "1010010110000" => data <= "000000";
				when "1010010110001" => data <= "000000";
				when "1010010110010" => data <= "000000";
				when "1010010110011" => data <= "111111";
				when "1010010110100" => data <= "100011";
				when "1010010110101" => data <= "100011";
				when "1010010110110" => data <= "111111";
				when "1010010110111" => data <= "000000";
				when "1010010111000" => data <= "000000";
				when "1010010111001" => data <= "000000";
				when "1010010111010" => data <= "000000";
				when "1010010111011" => data <= "000000";
				when "1010010111100" => data <= "000000";
				when "1010010111101" => data <= "000000";
				when "1010010111110" => data <= "000000";
				when "1010010111111" => data <= "111111";
				when "1010011000000" => data <= "100011";
				when "1010011000001" => data <= "100011";
				when "1010011000010" => data <= "111111";
				when "1010011000011" => data <= "000000";
				when "1010011000100" => data <= "000000";
				when "1010011000101" => data <= "000000";
				when "1010011000110" => data <= "000000";
				when "1010011000111" => data <= "111111";
				when "1010011001000" => data <= "100011";
				when "1010011001001" => data <= "100011";
				when "1010011001010" => data <= "111111";
				when "1010011001011" => data <= "000000";
				when "1010011001100" => data <= "000000";
				when "1010011001101" => data <= "000000";
				when "1010011001110" => data <= "000000";
				when "1010011001111" => data <= "000000";
				when "1010011010000" => data <= "000000";
				when "1010011010001" => data <= "000000";
				when "1010011010010" => data <= "000000";
				when "1010011010011" => data <= "111111";
				when "1010011010100" => data <= "100011";
				when "1010011010101" => data <= "100011";
				when "1010011010110" => data <= "111111";
				when "1010011010111" => data <= "000000";
				when "1010011011000" => data <= "000000";
				when "1010011011001" => data <= "000000";
				when "1010011011010" => data <= "000000";
				when "1010011011011" => data <= "000000";
				when "1010011011100" => data <= "000000";
				when "1010011011101" => data <= "000000";
				when "1010011011110" => data <= "000000";
				when "1010011011111" => data <= "000000";
				when "1010011100000" => data <= "000000";
				when "1010011100001" => data <= "111111";
				when "1010011100010" => data <= "100011";
				when "1010011100011" => data <= "100011";
				when "1010011100100" => data <= "111111";
				when "1010011100101" => data <= "000000";
				when "1010011100110" => data <= "000000";
				when "1010011100111" => data <= "000000";
				when "1010011101000" => data <= "000000";
				when "1010011101001" => data <= "111111";
				when "1010011101010" => data <= "100011";
				when "1010011101011" => data <= "100011";
				when "1010011101100" => data <= "111111";
				when "1010011101101" => data <= "000000";
				when "1010011101110" => data <= "000000";
				when "1010011101111" => data <= "000000";
				when "1010011110000" => data <= "000000";
				when "1010011110001" => data <= "000000";
				when "1010011110010" => data <= "000000";
				when "1010011110011" => data <= "000000";
				when "1010011110100" => data <= "000000";
				when "1010011110101" => data <= "000000";
				when "1010011110110" => data <= "000000";
				when "1010011110111" => data <= "000000";
				when "1010011111000" => data <= "000000";
				when "1010011111001" => data <= "000000";
				when "1010011111010" => data <= "000000";
				when "1010011111011" => data <= "000000";
				when "1010011111100" => data <= "000000";
				when "1010011111101" => data <= "000000";
				when "1010011111110" => data <= "000000";
				when "1010011111111" => data <= "000000";
				when "1010100000000" => data <= "000000";
				when "1010100000001" => data <= "000000";
				when "1010100000010" => data <= "000000";
				when "1010100000011" => data <= "000000";
				when "1010100000100" => data <= "000000";
				when "1010100000101" => data <= "000000";
				when "1010100000110" => data <= "000000";
				when "1010100000111" => data <= "000000";
				when "1010100001000" => data <= "000000";
				when "1010100001001" => data <= "000000";
				when "1010100001010" => data <= "000000";
				when "1010100001011" => data <= "000000";
				when "1010100001100" => data <= "000000";
				when "1010100001101" => data <= "111111";
				when "1010100001110" => data <= "100011";
				when "1010100001111" => data <= "100011";
				when "1010100010000" => data <= "111111";
				when "1010100010001" => data <= "000000";
				when "1010100010010" => data <= "000000";
				when "1010100010011" => data <= "000000";
				when "1010100010100" => data <= "000000";
				when "1010100010101" => data <= "111111";
				when "1010100010110" => data <= "100011";
				when "1010100010111" => data <= "100011";
				when "1010100011000" => data <= "111111";
				when "1010100011001" => data <= "000000";
				when "1010100011010" => data <= "000000";
				when "1010100011011" => data <= "000000";
				when "1010100011100" => data <= "000000";
				when "1010100011101" => data <= "000000";
				when "1010100011110" => data <= "000000";
				when "1010100011111" => data <= "000000";
				when "1010100100000" => data <= "000000";
				when "1010100100001" => data <= "000000";
				when "1010100100010" => data <= "111111";
				when "1010100100011" => data <= "100011";
				when "1010100100100" => data <= "100011";
				when "1010100100101" => data <= "111111";
				when "1010100100110" => data <= "000000";
				when "1010100100111" => data <= "000000";
				when "1010100101000" => data <= "000000";
				when "1010100101001" => data <= "000000";
				when "1010100101010" => data <= "000000";
				when "1010100101011" => data <= "000000";
				when "1010100101100" => data <= "000000";
				when "1010100101101" => data <= "000000";
				when "1010100101110" => data <= "000000";
				when "1010100101111" => data <= "000000";
				when "1010100110000" => data <= "000000";
				when "1010100110001" => data <= "000000";
				when "1010100110010" => data <= "000000";
				when "1010100110011" => data <= "111111";
				when "1010100110100" => data <= "100011";
				when "1010100110101" => data <= "100011";
				when "1010100110110" => data <= "111111";
				when "1010100110111" => data <= "000000";
				when "1010100111000" => data <= "000000";
				when "1010100111001" => data <= "000000";
				when "1010100111010" => data <= "000000";
				when "1010100111011" => data <= "000000";
				when "1010100111100" => data <= "000000";
				when "1010100111101" => data <= "000000";
				when "1010100111110" => data <= "000000";
				when "1010100111111" => data <= "111111";
				when "1010101000000" => data <= "100011";
				when "1010101000001" => data <= "100011";
				when "1010101000010" => data <= "111111";
				when "1010101000011" => data <= "000000";
				when "1010101000100" => data <= "000000";
				when "1010101000101" => data <= "000000";
				when "1010101000110" => data <= "000000";
				when "1010101000111" => data <= "111111";
				when "1010101001000" => data <= "100011";
				when "1010101001001" => data <= "100011";
				when "1010101001010" => data <= "111111";
				when "1010101001011" => data <= "000000";
				when "1010101001100" => data <= "000000";
				when "1010101001101" => data <= "000000";
				when "1010101001110" => data <= "000000";
				when "1010101001111" => data <= "000000";
				when "1010101010000" => data <= "000000";
				when "1010101010001" => data <= "000000";
				when "1010101010010" => data <= "000000";
				when "1010101010011" => data <= "111111";
				when "1010101010100" => data <= "100011";
				when "1010101010101" => data <= "100011";
				when "1010101010110" => data <= "111111";
				when "1010101010111" => data <= "000000";
				when "1010101011000" => data <= "000000";
				when "1010101011001" => data <= "000000";
				when "1010101011010" => data <= "000000";
				when "1010101011011" => data <= "000000";
				when "1010101011100" => data <= "000000";
				when "1010101011101" => data <= "000000";
				when "1010101011110" => data <= "000000";
				when "1010101011111" => data <= "000000";
				when "1010101100000" => data <= "000000";
				when "1010101100001" => data <= "111111";
				when "1010101100010" => data <= "100011";
				when "1010101100011" => data <= "100011";
				when "1010101100100" => data <= "111111";
				when "1010101100101" => data <= "000000";
				when "1010101100110" => data <= "000000";
				when "1010101100111" => data <= "000000";
				when "1010101101000" => data <= "000000";
				when "1010101101001" => data <= "111111";
				when "1010101101010" => data <= "100011";
				when "1010101101011" => data <= "100011";
				when "1010101101100" => data <= "111111";
				when "1010101101101" => data <= "000000";
				when "1010101101110" => data <= "000000";
				when "1010101101111" => data <= "000000";
				when "1010101110000" => data <= "000000";
				when "1010101110001" => data <= "000000";
				when "1010101110010" => data <= "000000";
				when "1010101110011" => data <= "000000";
				when "1010101110100" => data <= "000000";
				when "1010101110101" => data <= "000000";
				when "1010101110110" => data <= "000000";
				when "1010101110111" => data <= "000000";
				when "1010101111000" => data <= "000000";
				when "1010101111001" => data <= "000000";
				when "1010101111010" => data <= "000000";
				when "1010101111011" => data <= "000000";
				when "1010101111100" => data <= "000000";
				when "1010101111101" => data <= "000000";
				when "1010101111110" => data <= "000000";
				when "1010101111111" => data <= "000000";
				when "1010110000000" => data <= "000000";
				when "1010110000001" => data <= "000000";
				when "1010110000010" => data <= "000000";
				when "1010110000011" => data <= "000000";
				when "1010110000100" => data <= "000000";
				when "1010110000101" => data <= "000000";
				when "1010110000110" => data <= "000000";
				when "1010110000111" => data <= "000000";
				when "1010110001000" => data <= "000000";
				when "1010110001001" => data <= "000000";
				when "1010110001010" => data <= "000000";
				when "1010110001011" => data <= "000000";
				when "1010110001100" => data <= "000000";
				when "1010110001101" => data <= "111111";
				when "1010110001110" => data <= "100011";
				when "1010110001111" => data <= "100011";
				when "1010110010000" => data <= "111111";
				when "1010110010001" => data <= "000000";
				when "1010110010010" => data <= "000000";
				when "1010110010011" => data <= "000000";
				when "1010110010100" => data <= "000000";
				when "1010110010101" => data <= "111111";
				when "1010110010110" => data <= "100011";
				when "1010110010111" => data <= "100011";
				when "1010110011000" => data <= "111111";
				when "1010110011001" => data <= "000000";
				when "1010110011010" => data <= "000000";
				when "1010110011011" => data <= "000000";
				when "1010110011100" => data <= "000000";
				when "1010110011101" => data <= "000000";
				when "1010110011110" => data <= "000000";
				when "1010110011111" => data <= "000000";
				when "1010110100000" => data <= "000000";
				when "1010110100001" => data <= "000000";
				when "1010110100010" => data <= "111111";
				when "1010110100011" => data <= "100011";
				when "1010110100100" => data <= "100011";
				when "1010110100101" => data <= "111111";
				when "1010110100110" => data <= "000000";
				when "1010110100111" => data <= "000000";
				when "1010110101000" => data <= "000000";
				when "1010110101001" => data <= "000000";
				when "1010110101010" => data <= "000000";
				when "1010110101011" => data <= "000000";
				when "1010110101100" => data <= "000000";
				when "1010110101101" => data <= "000000";
				when "1010110101110" => data <= "000000";
				when "1010110101111" => data <= "000000";
				when "1010110110000" => data <= "000000";
				when "1010110110001" => data <= "000000";
				when "1010110110010" => data <= "000000";
				when "1010110110011" => data <= "111111";
				when "1010110110100" => data <= "100011";
				when "1010110110101" => data <= "100011";
				when "1010110110110" => data <= "111111";
				when "1010110110111" => data <= "000000";
				when "1010110111000" => data <= "000000";
				when "1010110111001" => data <= "000000";
				when "1010110111010" => data <= "000000";
				when "1010110111011" => data <= "000000";
				when "1010110111100" => data <= "000000";
				when "1010110111101" => data <= "000000";
				when "1010110111110" => data <= "000000";
				when "1010110111111" => data <= "111111";
				when "1010111000000" => data <= "100011";
				when "1010111000001" => data <= "100011";
				when "1010111000010" => data <= "111111";
				when "1010111000011" => data <= "000000";
				when "1010111000100" => data <= "000000";
				when "1010111000101" => data <= "000000";
				when "1010111000110" => data <= "000000";
				when "1010111000111" => data <= "111111";
				when "1010111001000" => data <= "100011";
				when "1010111001001" => data <= "100011";
				when "1010111001010" => data <= "111111";
				when "1010111001011" => data <= "000000";
				when "1010111001100" => data <= "000000";
				when "1010111001101" => data <= "000000";
				when "1010111001110" => data <= "000000";
				when "1010111001111" => data <= "000000";
				when "1010111010000" => data <= "000000";
				when "1010111010001" => data <= "000000";
				when "1010111010010" => data <= "000000";
				when "1010111010011" => data <= "111111";
				when "1010111010100" => data <= "100111";
				when "1010111010101" => data <= "100111";
				when "1010111010110" => data <= "111111";
				when "1010111010111" => data <= "000000";
				when "1010111011000" => data <= "000000";
				when "1010111011001" => data <= "000000";
				when "1010111011010" => data <= "000000";
				when "1010111011011" => data <= "000000";
				when "1010111011100" => data <= "000000";
				when "1010111011101" => data <= "000000";
				when "1010111011110" => data <= "000000";
				when "1010111011111" => data <= "000000";
				when "1010111100000" => data <= "000000";
				when "1010111100001" => data <= "111111";
				when "1010111100010" => data <= "100111";
				when "1010111100011" => data <= "100111";
				when "1010111100100" => data <= "111111";
				when "1010111100101" => data <= "000000";
				when "1010111100110" => data <= "000000";
				when "1010111100111" => data <= "000000";
				when "1010111101000" => data <= "000000";
				when "1010111101001" => data <= "111111";
				when "1010111101010" => data <= "100111";
				when "1010111101011" => data <= "100111";
				when "1010111101100" => data <= "111111";
				when "1010111101101" => data <= "000000";
				when "1010111101110" => data <= "000000";
				when "1010111101111" => data <= "000000";
				when "1010111110000" => data <= "000000";
				when "1010111110001" => data <= "000000";
				when "1010111110010" => data <= "000000";
				when "1010111110011" => data <= "000000";
				when "1010111110100" => data <= "000000";
				when "1010111110101" => data <= "000000";
				when "1010111110110" => data <= "000000";
				when "1010111110111" => data <= "000000";
				when "1010111111000" => data <= "000000";
				when "1010111111001" => data <= "000000";
				when "1010111111010" => data <= "000000";
				when "1010111111011" => data <= "000000";
				when "1010111111100" => data <= "000000";
				when "1010111111101" => data <= "000000";
				when "1010111111110" => data <= "000000";
				when "1010111111111" => data <= "000000";
				when "1011000000000" => data <= "000000";
				when "1011000000001" => data <= "000000";
				when "1011000000010" => data <= "000000";
				when "1011000000011" => data <= "000000";
				when "1011000000100" => data <= "000000";
				when "1011000000101" => data <= "000000";
				when "1011000000110" => data <= "000000";
				when "1011000000111" => data <= "000000";
				when "1011000001000" => data <= "000000";
				when "1011000001001" => data <= "000000";
				when "1011000001010" => data <= "000000";
				when "1011000001011" => data <= "000000";
				when "1011000001100" => data <= "000000";
				when "1011000001101" => data <= "111111";
				when "1011000001110" => data <= "100111";
				when "1011000001111" => data <= "100111";
				when "1011000010000" => data <= "111111";
				when "1011000010001" => data <= "000000";
				when "1011000010010" => data <= "000000";
				when "1011000010011" => data <= "000000";
				when "1011000010100" => data <= "000000";
				when "1011000010101" => data <= "111111";
				when "1011000010110" => data <= "100111";
				when "1011000010111" => data <= "100111";
				when "1011000011000" => data <= "111111";
				when "1011000011001" => data <= "000000";
				when "1011000011010" => data <= "000000";
				when "1011000011011" => data <= "000000";
				when "1011000011100" => data <= "000000";
				when "1011000011101" => data <= "000000";
				when "1011000011110" => data <= "000000";
				when "1011000011111" => data <= "000000";
				when "1011000100000" => data <= "000000";
				when "1011000100001" => data <= "000000";
				when "1011000100010" => data <= "111111";
				when "1011000100011" => data <= "100111";
				when "1011000100100" => data <= "100111";
				when "1011000100101" => data <= "111111";
				when "1011000100110" => data <= "000000";
				when "1011000100111" => data <= "000000";
				when "1011000101000" => data <= "000000";
				when "1011000101001" => data <= "000000";
				when "1011000101010" => data <= "000000";
				when "1011000101011" => data <= "000000";
				when "1011000101100" => data <= "000000";
				when "1011000101101" => data <= "000000";
				when "1011000101110" => data <= "000000";
				when "1011000101111" => data <= "000000";
				when "1011000110000" => data <= "000000";
				when "1011000110001" => data <= "000000";
				when "1011000110010" => data <= "000000";
				when "1011000110011" => data <= "111111";
				when "1011000110100" => data <= "100111";
				when "1011000110101" => data <= "100111";
				when "1011000110110" => data <= "111111";
				when "1011000110111" => data <= "000000";
				when "1011000111000" => data <= "000000";
				when "1011000111001" => data <= "000000";
				when "1011000111010" => data <= "000000";
				when "1011000111011" => data <= "000000";
				when "1011000111100" => data <= "000000";
				when "1011000111101" => data <= "000000";
				when "1011000111110" => data <= "000000";
				when "1011000111111" => data <= "111111";
				when "1011001000000" => data <= "100111";
				when "1011001000001" => data <= "100111";
				when "1011001000010" => data <= "111111";
				when "1011001000011" => data <= "000000";
				when "1011001000100" => data <= "000000";
				when "1011001000101" => data <= "000000";
				when "1011001000110" => data <= "000000";
				when "1011001000111" => data <= "111111";
				when "1011001001000" => data <= "100111";
				when "1011001001001" => data <= "100111";
				when "1011001001010" => data <= "111111";
				when "1011001001011" => data <= "000000";
				when "1011001001100" => data <= "000000";
				when "1011001001101" => data <= "000000";
				when "1011001001110" => data <= "000000";
				when "1011001001111" => data <= "000000";
				when "1011001010000" => data <= "000000";
				when "1011001010001" => data <= "000000";
				when "1011001010010" => data <= "000000";
				when "1011001010011" => data <= "111111";
				when "1011001010100" => data <= "100111";
				when "1011001010101" => data <= "100111";
				when "1011001010110" => data <= "111111";
				when "1011001010111" => data <= "000000";
				when "1011001011000" => data <= "000000";
				when "1011001011001" => data <= "000000";
				when "1011001011010" => data <= "000000";
				when "1011001011011" => data <= "000000";
				when "1011001011100" => data <= "000000";
				when "1011001011101" => data <= "000000";
				when "1011001011110" => data <= "000000";
				when "1011001011111" => data <= "000000";
				when "1011001100000" => data <= "000000";
				when "1011001100001" => data <= "111111";
				when "1011001100010" => data <= "100111";
				when "1011001100011" => data <= "100111";
				when "1011001100100" => data <= "111111";
				when "1011001100101" => data <= "000000";
				when "1011001100110" => data <= "000000";
				when "1011001100111" => data <= "000000";
				when "1011001101000" => data <= "000000";
				when "1011001101001" => data <= "111111";
				when "1011001101010" => data <= "100111";
				when "1011001101011" => data <= "100111";
				when "1011001101100" => data <= "111111";
				when "1011001101101" => data <= "000000";
				when "1011001101110" => data <= "000000";
				when "1011001101111" => data <= "000000";
				when "1011001110000" => data <= "000000";
				when "1011001110001" => data <= "000000";
				when "1011001110010" => data <= "000000";
				when "1011001110011" => data <= "000000";
				when "1011001110100" => data <= "000000";
				when "1011001110101" => data <= "000000";
				when "1011001110110" => data <= "000000";
				when "1011001110111" => data <= "000000";
				when "1011001111000" => data <= "000000";
				when "1011001111001" => data <= "000000";
				when "1011001111010" => data <= "000000";
				when "1011001111011" => data <= "000000";
				when "1011001111100" => data <= "000000";
				when "1011001111101" => data <= "000000";
				when "1011001111110" => data <= "000000";
				when "1011001111111" => data <= "000000";
				when "1011010000000" => data <= "000000";
				when "1011010000001" => data <= "000000";
				when "1011010000010" => data <= "000000";
				when "1011010000011" => data <= "000000";
				when "1011010000100" => data <= "000000";
				when "1011010000101" => data <= "000000";
				when "1011010000110" => data <= "000000";
				when "1011010000111" => data <= "000000";
				when "1011010001000" => data <= "000000";
				when "1011010001001" => data <= "000000";
				when "1011010001010" => data <= "000000";
				when "1011010001011" => data <= "000000";
				when "1011010001100" => data <= "000000";
				when "1011010001101" => data <= "111111";
				when "1011010001110" => data <= "100111";
				when "1011010001111" => data <= "100111";
				when "1011010010000" => data <= "111111";
				when "1011010010001" => data <= "000000";
				when "1011010010010" => data <= "000000";
				when "1011010010011" => data <= "000000";
				when "1011010010100" => data <= "000000";
				when "1011010010101" => data <= "111111";
				when "1011010010110" => data <= "100111";
				when "1011010010111" => data <= "100111";
				when "1011010011000" => data <= "111111";
				when "1011010011001" => data <= "000000";
				when "1011010011010" => data <= "000000";
				when "1011010011011" => data <= "000000";
				when "1011010011100" => data <= "000000";
				when "1011010011101" => data <= "000000";
				when "1011010011110" => data <= "000000";
				when "1011010011111" => data <= "000000";
				when "1011010100000" => data <= "000000";
				when "1011010100001" => data <= "000000";
				when "1011010100010" => data <= "111111";
				when "1011010100011" => data <= "100111";
				when "1011010100100" => data <= "100111";
				when "1011010100101" => data <= "111111";
				when "1011010100110" => data <= "000000";
				when "1011010100111" => data <= "000000";
				when "1011010101000" => data <= "000000";
				when "1011010101001" => data <= "000000";
				when "1011010101010" => data <= "000000";
				when "1011010101011" => data <= "000000";
				when "1011010101100" => data <= "000000";
				when "1011010101101" => data <= "000000";
				when "1011010101110" => data <= "000000";
				when "1011010101111" => data <= "000000";
				when "1011010110000" => data <= "000000";
				when "1011010110001" => data <= "000000";
				when "1011010110010" => data <= "000000";
				when "1011010110011" => data <= "111111";
				when "1011010110100" => data <= "100111";
				when "1011010110101" => data <= "100111";
				when "1011010110110" => data <= "111111";
				when "1011010110111" => data <= "000000";
				when "1011010111000" => data <= "000000";
				when "1011010111001" => data <= "000000";
				when "1011010111010" => data <= "000000";
				when "1011010111011" => data <= "000000";
				when "1011010111100" => data <= "000000";
				when "1011010111101" => data <= "000000";
				when "1011010111110" => data <= "000000";
				when "1011010111111" => data <= "111111";
				when "1011011000000" => data <= "100111";
				when "1011011000001" => data <= "100111";
				when "1011011000010" => data <= "111111";
				when "1011011000011" => data <= "000000";
				when "1011011000100" => data <= "000000";
				when "1011011000101" => data <= "000000";
				when "1011011000110" => data <= "000000";
				when "1011011000111" => data <= "111111";
				when "1011011001000" => data <= "100111";
				when "1011011001001" => data <= "100111";
				when "1011011001010" => data <= "111111";
				when "1011011001011" => data <= "000000";
				when "1011011001100" => data <= "000000";
				when "1011011001101" => data <= "000000";
				when "1011011001110" => data <= "000000";
				when "1011011001111" => data <= "000000";
				when "1011011010000" => data <= "000000";
				when "1011011010001" => data <= "000000";
				when "1011011010010" => data <= "000000";
				when "1011011010011" => data <= "111111";
				when "1011011010100" => data <= "100111";
				when "1011011010101" => data <= "100111";
				when "1011011010110" => data <= "111111";
				when "1011011010111" => data <= "000000";
				when "1011011011000" => data <= "000000";
				when "1011011011001" => data <= "000000";
				when "1011011011010" => data <= "000000";
				when "1011011011011" => data <= "000000";
				when "1011011011100" => data <= "000000";
				when "1011011011101" => data <= "000000";
				when "1011011011110" => data <= "000000";
				when "1011011011111" => data <= "000000";
				when "1011011100000" => data <= "000000";
				when "1011011100001" => data <= "111111";
				when "1011011100010" => data <= "100111";
				when "1011011100011" => data <= "100111";
				when "1011011100100" => data <= "111111";
				when "1011011100101" => data <= "000000";
				when "1011011100110" => data <= "000000";
				when "1011011100111" => data <= "000000";
				when "1011011101000" => data <= "000000";
				when "1011011101001" => data <= "111111";
				when "1011011101010" => data <= "100111";
				when "1011011101011" => data <= "100111";
				when "1011011101100" => data <= "111111";
				when "1011011101101" => data <= "000000";
				when "1011011101110" => data <= "000000";
				when "1011011101111" => data <= "000000";
				when "1011011110000" => data <= "000000";
				when "1011011110001" => data <= "000000";
				when "1011011110010" => data <= "000000";
				when "1011011110011" => data <= "000000";
				when "1011011110100" => data <= "000000";
				when "1011011110101" => data <= "000000";
				when "1011011110110" => data <= "000000";
				when "1011011110111" => data <= "000000";
				when "1011011111000" => data <= "000000";
				when "1011011111001" => data <= "000000";
				when "1011011111010" => data <= "000000";
				when "1011011111011" => data <= "000000";
				when "1011011111100" => data <= "000000";
				when "1011011111101" => data <= "000000";
				when "1011011111110" => data <= "000000";
				when "1011011111111" => data <= "000000";
				when "1011100000000" => data <= "000000";
				when "1011100000001" => data <= "000000";
				when "1011100000010" => data <= "000000";
				when "1011100000011" => data <= "000000";
				when "1011100000100" => data <= "000000";
				when "1011100000101" => data <= "000000";
				when "1011100000110" => data <= "000000";
				when "1011100000111" => data <= "000000";
				when "1011100001000" => data <= "000000";
				when "1011100001001" => data <= "000000";
				when "1011100001010" => data <= "000000";
				when "1011100001011" => data <= "000000";
				when "1011100001100" => data <= "000000";
				when "1011100001101" => data <= "111111";
				when "1011100001110" => data <= "100111";
				when "1011100001111" => data <= "100111";
				when "1011100010000" => data <= "111111";
				when "1011100010001" => data <= "000000";
				when "1011100010010" => data <= "000000";
				when "1011100010011" => data <= "000000";
				when "1011100010100" => data <= "000000";
				when "1011100010101" => data <= "111111";
				when "1011100010110" => data <= "100111";
				when "1011100010111" => data <= "100111";
				when "1011100011000" => data <= "111111";
				when "1011100011001" => data <= "000000";
				when "1011100011010" => data <= "000000";
				when "1011100011011" => data <= "000000";
				when "1011100011100" => data <= "000000";
				when "1011100011101" => data <= "000000";
				when "1011100011110" => data <= "000000";
				when "1011100011111" => data <= "000000";
				when "1011100100000" => data <= "000000";
				when "1011100100001" => data <= "000000";
				when "1011100100010" => data <= "111111";
				when "1011100100011" => data <= "100111";
				when "1011100100100" => data <= "100111";
				when "1011100100101" => data <= "111111";
				when "1011100100110" => data <= "000000";
				when "1011100100111" => data <= "000000";
				when "1011100101000" => data <= "000000";
				when "1011100101001" => data <= "000000";
				when "1011100101010" => data <= "000000";
				when "1011100101011" => data <= "000000";
				when "1011100101100" => data <= "000000";
				when "1011100101101" => data <= "000000";
				when "1011100101110" => data <= "000000";
				when "1011100101111" => data <= "000000";
				when "1011100110000" => data <= "000000";
				when "1011100110001" => data <= "000000";
				when "1011100110010" => data <= "000000";
				when "1011100110011" => data <= "111111";
				when "1011100110100" => data <= "100111";
				when "1011100110101" => data <= "100111";
				when "1011100110110" => data <= "111111";
				when "1011100110111" => data <= "000000";
				when "1011100111000" => data <= "000000";
				when "1011100111001" => data <= "000000";
				when "1011100111010" => data <= "000000";
				when "1011100111011" => data <= "000000";
				when "1011100111100" => data <= "000000";
				when "1011100111101" => data <= "000000";
				when "1011100111110" => data <= "000000";
				when "1011100111111" => data <= "111111";
				when "1011101000000" => data <= "100111";
				when "1011101000001" => data <= "100111";
				when "1011101000010" => data <= "111111";
				when "1011101000011" => data <= "000000";
				when "1011101000100" => data <= "000000";
				when "1011101000101" => data <= "000000";
				when "1011101000110" => data <= "000000";
				when "1011101000111" => data <= "111111";
				when "1011101001000" => data <= "100111";
				when "1011101001001" => data <= "100111";
				when "1011101001010" => data <= "111111";
				when "1011101001011" => data <= "000000";
				when "1011101001100" => data <= "000000";
				when "1011101001101" => data <= "000000";
				when "1011101001110" => data <= "000000";
				when "1011101001111" => data <= "000000";
				when "1011101010000" => data <= "000000";
				when "1011101010001" => data <= "000000";
				when "1011101010010" => data <= "000000";
				when "1011101010011" => data <= "000000";
				when "1011101010100" => data <= "111111";
				when "1011101010101" => data <= "111111";
				when "1011101010110" => data <= "000000";
				when "1011101010111" => data <= "000000";
				when "1011101011000" => data <= "000000";
				when "1011101011001" => data <= "000000";
				when "1011101011010" => data <= "000000";
				when "1011101011011" => data <= "000000";
				when "1011101011100" => data <= "000000";
				when "1011101011101" => data <= "000000";
				when "1011101011110" => data <= "000000";
				when "1011101011111" => data <= "000000";
				when "1011101100000" => data <= "000000";
				when "1011101100001" => data <= "000000";
				when "1011101100010" => data <= "111111";
				when "1011101100011" => data <= "111111";
				when "1011101100100" => data <= "000000";
				when "1011101100101" => data <= "000000";
				when "1011101100110" => data <= "000000";
				when "1011101100111" => data <= "000000";
				when "1011101101000" => data <= "000000";
				when "1011101101001" => data <= "000000";
				when "1011101101010" => data <= "111111";
				when "1011101101011" => data <= "111111";
				when "1011101101100" => data <= "000000";
				when "1011101101101" => data <= "000000";
				when "1011101101110" => data <= "000000";
				when "1011101101111" => data <= "000000";
				when "1011101110000" => data <= "000000";
				when "1011101110001" => data <= "000000";
				when "1011101110010" => data <= "000000";
				when "1011101110011" => data <= "000000";
				when "1011101110100" => data <= "000000";
				when "1011101110101" => data <= "000000";
				when "1011101110110" => data <= "000000";
				when "1011101110111" => data <= "000000";
				when "1011101111000" => data <= "000000";
				when "1011101111001" => data <= "000000";
				when "1011101111010" => data <= "000000";
				when "1011101111011" => data <= "000000";
				when "1011101111100" => data <= "000000";
				when "1011101111101" => data <= "000000";
				when "1011101111110" => data <= "000000";
				when "1011101111111" => data <= "000000";
				when "1011110000000" => data <= "000000";
				when "1011110000001" => data <= "000000";
				when "1011110000010" => data <= "000000";
				when "1011110000011" => data <= "000000";
				when "1011110000100" => data <= "000000";
				when "1011110000101" => data <= "000000";
				when "1011110000110" => data <= "000000";
				when "1011110000111" => data <= "000000";
				when "1011110001000" => data <= "000000";
				when "1011110001001" => data <= "000000";
				when "1011110001010" => data <= "000000";
				when "1011110001011" => data <= "000000";
				when "1011110001100" => data <= "000000";
				when "1011110001101" => data <= "000000";
				when "1011110001110" => data <= "111111";
				when "1011110001111" => data <= "111111";
				when "1011110010000" => data <= "000000";
				when "1011110010001" => data <= "000000";
				when "1011110010010" => data <= "000000";
				when "1011110010011" => data <= "000000";
				when "1011110010100" => data <= "000000";
				when "1011110010101" => data <= "000000";
				when "1011110010110" => data <= "111111";
				when "1011110010111" => data <= "111111";
				when "1011110011000" => data <= "000000";
				when "1011110011001" => data <= "000000";
				when "1011110011010" => data <= "000000";
				when "1011110011011" => data <= "000000";
				when "1011110011100" => data <= "000000";
				when "1011110011101" => data <= "000000";
				when "1011110011110" => data <= "000000";
				when "1011110011111" => data <= "000000";
				when "1011110100000" => data <= "000000";
				when "1011110100001" => data <= "000000";
				when "1011110100010" => data <= "000000";
				when "1011110100011" => data <= "111111";
				when "1011110100100" => data <= "111111";
				when "1011110100101" => data <= "000000";
				when "1011110100110" => data <= "000000";
				when "1011110100111" => data <= "000000";
				when "1011110101000" => data <= "000000";
				when "1011110101001" => data <= "000000";
				when "1011110101010" => data <= "000000";
				when "1011110101011" => data <= "000000";
				when "1011110101100" => data <= "000000";
				when "1011110101101" => data <= "000000";
				when "1011110101110" => data <= "000000";
				when "1011110101111" => data <= "000000";
				when "1011110110000" => data <= "000000";
				when "1011110110001" => data <= "000000";
				when "1011110110010" => data <= "000000";
				when "1011110110011" => data <= "000000";
				when "1011110110100" => data <= "111111";
				when "1011110110101" => data <= "111111";
				when "1011110110110" => data <= "000000";
				when "1011110110111" => data <= "000000";
				when "1011110111000" => data <= "000000";
				when "1011110111001" => data <= "000000";
				when "1011110111010" => data <= "000000";
				when "1011110111011" => data <= "000000";
				when "1011110111100" => data <= "000000";
				when "1011110111101" => data <= "000000";
				when "1011110111110" => data <= "000000";
				when "1011110111111" => data <= "000000";
				when "1011111000000" => data <= "111111";
				when "1011111000001" => data <= "111111";
				when "1011111000010" => data <= "000000";
				when "1011111000011" => data <= "000000";
				when "1011111000100" => data <= "000000";
				when "1011111000101" => data <= "000000";
				when "1011111000110" => data <= "000000";
				when "1011111000111" => data <= "000000";
				when "1011111001000" => data <= "111111";
				when "1011111001001" => data <= "111111";
				when "1011111001010" => data <= "000000";
				when "1011111001011" => data <= "000000";
				when "1011111001100" => data <= "000000";
				when "1011111001101" => data <= "000000";
				when "1011111001110" => data <= "000000";
				when "1011111001111" => data <= "000000";
				when "1011111010000" => data <= "000000";
				when "1011111010001" => data <= "000000";
				when "1011111010010" => data <= "000000";
				when "1011111010011" => data <= "000000";
				when "1011111010100" => data <= "000000";
				when "1011111010101" => data <= "000000";
				when "1011111010110" => data <= "000000";
				when "1011111010111" => data <= "000000";
				when "1011111011000" => data <= "000000";
				when "1011111011001" => data <= "000000";
				when "1011111011010" => data <= "000000";
				when "1011111011011" => data <= "000000";
				when "1011111011100" => data <= "000000";
				when "1011111011101" => data <= "000000";
				when "1011111011110" => data <= "000000";
				when "1011111011111" => data <= "000000";
				when "1011111100000" => data <= "000000";
				when "1011111100001" => data <= "000000";
				when "1011111100010" => data <= "000000";
				when "1011111100011" => data <= "000000";
				when "1011111100100" => data <= "000000";
				when "1011111100101" => data <= "000000";
				when "1011111100110" => data <= "000000";
				when "1011111100111" => data <= "000000";
				when "1011111101000" => data <= "000000";
				when "1011111101001" => data <= "000000";
				when "1011111101010" => data <= "000000";
				when "1011111101011" => data <= "000000";
				when "1011111101100" => data <= "000000";
				when "1011111101101" => data <= "000000";
				when "1011111101110" => data <= "000000";
				when "1011111101111" => data <= "000000";
				when "1011111110000" => data <= "000000";
				when "1011111110001" => data <= "000000";
				when "1011111110010" => data <= "000000";
				when "1011111110011" => data <= "000000";
				when "1011111110100" => data <= "000000";
				when "1011111110101" => data <= "000000";
				when "1011111110110" => data <= "000000";
				when "1011111110111" => data <= "000000";
				when "1011111111000" => data <= "000000";
				when "1011111111001" => data <= "000000";
				when "1011111111010" => data <= "000000";
				when "1011111111011" => data <= "000000";
				when "1011111111100" => data <= "000000";
				when "1011111111101" => data <= "000000";
				when "1011111111110" => data <= "000000";
				when "1011111111111" => data <= "000000";
				when "1100000000000" => data <= "000000";
				when "1100000000001" => data <= "000000";
				when "1100000000010" => data <= "000000";
				when "1100000000011" => data <= "000000";
				when "1100000000100" => data <= "000000";
				when "1100000000101" => data <= "000000";
				when "1100000000110" => data <= "000000";
				when "1100000000111" => data <= "000000";
				when "1100000001000" => data <= "000000";
				when "1100000001001" => data <= "000000";
				when "1100000001010" => data <= "000000";
				when "1100000001011" => data <= "000000";
				when "1100000001100" => data <= "000000";
				when "1100000001101" => data <= "000000";
				when "1100000001110" => data <= "000000";
				when "1100000001111" => data <= "000000";
				when "1100000010000" => data <= "000000";
				when "1100000010001" => data <= "000000";
				when "1100000010010" => data <= "000000";
				when "1100000010011" => data <= "000000";
				when "1100000010100" => data <= "000000";
				when "1100000010101" => data <= "000000";
				when "1100000010110" => data <= "000000";
				when "1100000010111" => data <= "000000";
				when "1100000011000" => data <= "000000";
				when "1100000011001" => data <= "000000";
				when "1100000011010" => data <= "000000";
				when "1100000011011" => data <= "000000";
				when "1100000011100" => data <= "000000";
				when "1100000011101" => data <= "000000";
				when "1100000011110" => data <= "000000";
				when "1100000011111" => data <= "000000";
				when "1100000100000" => data <= "000000";
				when "1100000100001" => data <= "000000";
				when "1100000100010" => data <= "000000";
				when "1100000100011" => data <= "000000";
				when "1100000100100" => data <= "000000";
				when "1100000100101" => data <= "000000";
				when "1100000100110" => data <= "000000";
				when "1100000100111" => data <= "000000";
				when "1100000101000" => data <= "000000";
				when "1100000101001" => data <= "000000";
				when "1100000101010" => data <= "000000";
				when "1100000101011" => data <= "000000";
				when "1100000101100" => data <= "000000";
				when "1100000101101" => data <= "000000";
				when "1100000101110" => data <= "000000";
				when "1100000101111" => data <= "000000";
				when "1100000110000" => data <= "000000";
				when "1100000110001" => data <= "000000";
				when "1100000110010" => data <= "000000";
				when "1100000110011" => data <= "000000";
				when "1100000110100" => data <= "000000";
				when "1100000110101" => data <= "000000";
				when "1100000110110" => data <= "000000";
				when "1100000110111" => data <= "000000";
				when "1100000111000" => data <= "000000";
				when "1100000111001" => data <= "000000";
				when "1100000111010" => data <= "000000";
				when "1100000111011" => data <= "000000";
				when "1100000111100" => data <= "000000";
				when "1100000111101" => data <= "000000";
				when "1100000111110" => data <= "000000";
				when "1100000111111" => data <= "000000";
				when "1100001000000" => data <= "000000";
				when "1100001000001" => data <= "000000";
				when "1100001000010" => data <= "000000";
				when "1100001000011" => data <= "000000";
				when "1100001000100" => data <= "000000";
				when "1100001000101" => data <= "000000";
				when "1100001000110" => data <= "000000";
				when "1100001000111" => data <= "000000";
				when "1100001001000" => data <= "000000";
				when "1100001001001" => data <= "000000";
				when "1100001001010" => data <= "000000";
				when "1100001001011" => data <= "000000";
				when "1100001001100" => data <= "000000";
				when "1100001001101" => data <= "000000";
				when "1100001001110" => data <= "000000";
				when "1100001001111" => data <= "000000";
				when "1100001010000" => data <= "000000";
				when "1100001010001" => data <= "000000";
				when "1100001010010" => data <= "000000";
				when "1100001010011" => data <= "000000";
				when "1100001010100" => data <= "000000";
				when "1100001010101" => data <= "000000";
				when "1100001010110" => data <= "000000";
				when "1100001010111" => data <= "000000";
				when "1100001011000" => data <= "000000";
				when "1100001011001" => data <= "000000";
				when "1100001011010" => data <= "000000";
				when "1100001011011" => data <= "000000";
				when "1100001011100" => data <= "000000";
				when "1100001011101" => data <= "000000";
				when "1100001011110" => data <= "000000";
				when "1100001011111" => data <= "000000";
				when "1100001100000" => data <= "000000";
				when "1100001100001" => data <= "000000";
				when "1100001100010" => data <= "000000";
				when "1100001100011" => data <= "000000";
				when "1100001100100" => data <= "000000";
				when "1100001100101" => data <= "000000";
				when "1100001100110" => data <= "000000";
				when "1100001100111" => data <= "000000";
				when "1100001101000" => data <= "000000";
				when "1100001101001" => data <= "000000";
				when "1100001101010" => data <= "000000";
				when "1100001101011" => data <= "000000";
				when "1100001101100" => data <= "000000";
				when "1100001101101" => data <= "000000";
				when "1100001101110" => data <= "000000";
				when "1100001101111" => data <= "000000";
				when "1100001110000" => data <= "000000";
				when "1100001110001" => data <= "000000";
				when "1100001110010" => data <= "000000";
				when "1100001110011" => data <= "000000";
				when "1100001110100" => data <= "000000";
				when "1100001110101" => data <= "000000";
				when "1100001110110" => data <= "000000";
				when "1100001110111" => data <= "000000";
				when "1100001111000" => data <= "000000";
				when "1100001111001" => data <= "000000";
				when "1100001111010" => data <= "000000";
				when "1100001111011" => data <= "000000";
				when "1100001111100" => data <= "000000";
				when "1100001111101" => data <= "000000";
				when "1100001111110" => data <= "000000";
				when "1100001111111" => data <= "000000";
				when "1100010000000" => data <= "000000";
				when "1100010000001" => data <= "000000";
				when "1100010000010" => data <= "000000";
				when "1100010000011" => data <= "000000";
				when "1100010000100" => data <= "000000";
				when "1100010000101" => data <= "000000";
				when "1100010000110" => data <= "000000";
				when "1100010000111" => data <= "000000";
				when "1100010001000" => data <= "000000";
				when "1100010001001" => data <= "000000";
				when "1100010001010" => data <= "000000";
				when "1100010001011" => data <= "000000";
				when "1100010001100" => data <= "000000";
				when "1100010001101" => data <= "000000";
				when "1100010001110" => data <= "000000";
				when "1100010001111" => data <= "000000";
				when "1100010010000" => data <= "000000";
				when "1100010010001" => data <= "000000";
				when "1100010010010" => data <= "000000";
				when "1100010010011" => data <= "000000";
				when "1100010010100" => data <= "000000";
				when "1100010010101" => data <= "000000";
				when "1100010010110" => data <= "000000";
				when "1100010010111" => data <= "000000";
				when "1100010011000" => data <= "000000";
				when "1100010011001" => data <= "000000";
				when "1100010011010" => data <= "000000";
				when "1100010011011" => data <= "000000";
				when "1100010011100" => data <= "000000";
				when "1100010011101" => data <= "000000";
				when "1100010011110" => data <= "000000";
				when "1100010011111" => data <= "000000";
				when "1100010100000" => data <= "000000";
				when "1100010100001" => data <= "000000";
				when "1100010100010" => data <= "000000";
				when "1100010100011" => data <= "000000";
				when "1100010100100" => data <= "000000";
				when "1100010100101" => data <= "000000";
				when "1100010100110" => data <= "000000";
				when "1100010100111" => data <= "000000";
				when "1100010101000" => data <= "000000";
				when "1100010101001" => data <= "000000";
				when "1100010101010" => data <= "000000";
				when "1100010101011" => data <= "000000";
				when "1100010101100" => data <= "000000";
				when "1100010101101" => data <= "000000";
				when "1100010101110" => data <= "000000";
				when "1100010101111" => data <= "000000";
				when "1100010110000" => data <= "000000";
				when "1100010110001" => data <= "000000";
				when "1100010110010" => data <= "000000";
				when "1100010110011" => data <= "000000";
				when "1100010110100" => data <= "000000";
				when "1100010110101" => data <= "000000";
				when "1100010110110" => data <= "000000";
				when "1100010110111" => data <= "000000";
				when "1100010111000" => data <= "000000";
				when "1100010111001" => data <= "000000";
				when "1100010111010" => data <= "000000";
				when "1100010111011" => data <= "000000";
				when "1100010111100" => data <= "000000";
				when "1100010111101" => data <= "000000";
				when "1100010111110" => data <= "000000";
				when "1100010111111" => data <= "000000";
				when "1100011000000" => data <= "000000";
				when "1100011000001" => data <= "000000";
				when "1100011000010" => data <= "000000";
				when "1100011000011" => data <= "000000";
				when "1100011000100" => data <= "000000";
				when "1100011000101" => data <= "000000";
				when "1100011000110" => data <= "000000";
				when "1100011000111" => data <= "000000";
				when "1100011001000" => data <= "000000";
				when "1100011001001" => data <= "000000";
				when "1100011001010" => data <= "000000";
				when "1100011001011" => data <= "000000";
				when "1100011001100" => data <= "000000";
				when "1100011001101" => data <= "000000";
				when "1100011001110" => data <= "000000";
				when "1100011001111" => data <= "000000";
				when "1100011010000" => data <= "000000";
				when "1100011010001" => data <= "010011";
				when "1100011010010" => data <= "000000";
				when "1100011010011" => data <= "000000";
				when "1100011010100" => data <= "000000";
				when "1100011010101" => data <= "000000";
				when "1100011010110" => data <= "000000";
				when "1100011010111" => data <= "000000";
				when "1100011011000" => data <= "000000";
				when "1100011011001" => data <= "000000";
				when "1100011011010" => data <= "000000";
				when "1100011011011" => data <= "000000";
				when "1100011011100" => data <= "000000";
				when "1100011011101" => data <= "000000";
				when "1100011011110" => data <= "000000";
				when "1100011011111" => data <= "000000";
				when "1100011100000" => data <= "000000";
				when "1100011100001" => data <= "000000";
				when "1100011100010" => data <= "000000";
				when "1100011100011" => data <= "000000";
				when "1100011100100" => data <= "000000";
				when "1100011100101" => data <= "000000";
				when "1100011100110" => data <= "000000";
				when "1100011100111" => data <= "000000";
				when "1100011101000" => data <= "000000";
				when "1100011101001" => data <= "000000";
				when "1100011101010" => data <= "000000";
				when "1100011101011" => data <= "000000";
				when "1100011101100" => data <= "000000";
				when "1100011101101" => data <= "000000";
				when "1100011101110" => data <= "000000";
				when "1100011101111" => data <= "000000";
				when "1100011110000" => data <= "000000";
				when "1100011110001" => data <= "000000";
				when "1100011110010" => data <= "000000";
				when "1100011110011" => data <= "000000";
				when "1100011110100" => data <= "000000";
				when "1100011110101" => data <= "000000";
				when "1100011110110" => data <= "000000";
				when "1100011110111" => data <= "000000";
				when "1100011111000" => data <= "000000";
				when "1100011111001" => data <= "000000";
				when "1100011111010" => data <= "000000";
				when "1100011111011" => data <= "000000";
				when "1100011111100" => data <= "000000";
				when "1100011111101" => data <= "000000";
				when "1100011111110" => data <= "000000";
				when "1100011111111" => data <= "000000";
				when "1100100000000" => data <= "000000";
				when "1100100000001" => data <= "000000";
				when "1100100000010" => data <= "000000";
				when "1100100000011" => data <= "000000";
				when "1100100000100" => data <= "000000";
				when "1100100000101" => data <= "000000";
				when "1100100000110" => data <= "000000";
				when "1100100000111" => data <= "000000";
				when "1100100001000" => data <= "000000";
				when "1100100001001" => data <= "000000";
				when "1100100001010" => data <= "000000";
				when "1100100001011" => data <= "000000";
				when "1100100001100" => data <= "000000";
				when "1100100001101" => data <= "000000";
				when "1100100001110" => data <= "000000";
				when "1100100001111" => data <= "000000";
				when "1100100010000" => data <= "000000";
				when "1100100010001" => data <= "000000";
				when "1100100010010" => data <= "000000";
				when "1100100010011" => data <= "000000";
				when "1100100010100" => data <= "000000";
				when "1100100010101" => data <= "000000";
				when "1100100010110" => data <= "000000";
				when "1100100010111" => data <= "000000";
				when "1100100011000" => data <= "000000";
				when "1100100011001" => data <= "000000";
				when "1100100011010" => data <= "000000";
				when "1100100011011" => data <= "000000";
				when "1100100011100" => data <= "000000";
				when "1100100011101" => data <= "000000";
				when "1100100011110" => data <= "000000";
				when "1100100011111" => data <= "000000";
				when "1100100100000" => data <= "000000";
				when "1100100100001" => data <= "000000";
				when "1100100100010" => data <= "000000";
				when "1100100100011" => data <= "000000";
				when "1100100100100" => data <= "000000";
				when "1100100100101" => data <= "000000";
				when "1100100100110" => data <= "000000";
				when "1100100100111" => data <= "000000";
				when "1100100101000" => data <= "000000";
				when "1100100101001" => data <= "000000";
				when "1100100101010" => data <= "000000";
				when "1100100101011" => data <= "000000";
				when "1100100101100" => data <= "000000";
				when "1100100101101" => data <= "000000";
				when "1100100101110" => data <= "000000";
				when "1100100101111" => data <= "010011";
				when "1100100110000" => data <= "010011";
				when "1100100110001" => data <= "010011";
				when "1100100110010" => data <= "010011";
				when "1100100110011" => data <= "010011";
				when "1100100110100" => data <= "000000";
				when "1100100110101" => data <= "000000";
				when "1100100110110" => data <= "000000";
				when "1100100110111" => data <= "000000";
				when "1100100111000" => data <= "000000";
				when "1100100111001" => data <= "000000";
				when "1100100111010" => data <= "000000";
				when "1100100111011" => data <= "000000";
				when "1100100111100" => data <= "000000";
				when "1100100111101" => data <= "000000";
				when "1100100111110" => data <= "000000";
				when "1100100111111" => data <= "000000";
				when "1100101000000" => data <= "000000";
				when "1100101000001" => data <= "000000";
				when "1100101000010" => data <= "000000";
				when "1100101000011" => data <= "000000";
				when "1100101000100" => data <= "000000";
				when "1100101000101" => data <= "000000";
				when "1100101000110" => data <= "000000";
				when "1100101000111" => data <= "000000";
				when "1100101001000" => data <= "000000";
				when "1100101001001" => data <= "000000";
				when "1100101001010" => data <= "000000";
				when "1100101001011" => data <= "000000";
				when "1100101001100" => data <= "000000";
				when "1100101001101" => data <= "000000";
				when "1100101001110" => data <= "000000";
				when "1100101001111" => data <= "000000";
				when "1100101010000" => data <= "000000";
				when "1100101010001" => data <= "010011";
				when "1100101010010" => data <= "000000";
				when "1100101010011" => data <= "000000";
				when "1100101010100" => data <= "000000";
				when "1100101010101" => data <= "000000";
				when "1100101010110" => data <= "000000";
				when "1100101010111" => data <= "000000";
				when "1100101011000" => data <= "000000";
				when "1100101011001" => data <= "000000";
				when "1100101011010" => data <= "000000";
				when "1100101011011" => data <= "000000";
				when "1100101011100" => data <= "000000";
				when "1100101011101" => data <= "000000";
				when "1100101011110" => data <= "000000";
				when "1100101011111" => data <= "000000";
				when "1100101100000" => data <= "000000";
				when "1100101100001" => data <= "000000";
				when "1100101100010" => data <= "000000";
				when "1100101100011" => data <= "000000";
				when "1100101100100" => data <= "000000";
				when "1100101100101" => data <= "000000";
				when "1100101100110" => data <= "000000";
				when "1100101100111" => data <= "000000";
				when "1100101101000" => data <= "000000";
				when "1100101101001" => data <= "000000";
				when "1100101101010" => data <= "000000";
				when "1100101101011" => data <= "000000";
				when "1100101101100" => data <= "000000";
				when "1100101101101" => data <= "000000";
				when "1100101101110" => data <= "000000";
				when "1100101101111" => data <= "000000";
				when "1100101110000" => data <= "000000";
				when "1100101110001" => data <= "000000";
				when "1100101110010" => data <= "000000";
				when "1100101110011" => data <= "000000";
				when "1100101110100" => data <= "000000";
				when "1100101110101" => data <= "000000";
				when "1100101110110" => data <= "000000";
				when "1100101110111" => data <= "000000";
				when "1100101111000" => data <= "000000";
				when "1100101111001" => data <= "000000";
				when "1100101111010" => data <= "000000";
				when "1100101111011" => data <= "000000";
				when "1100101111100" => data <= "000000";
				when "1100101111101" => data <= "000000";
				when "1100101111110" => data <= "000000";
				when "1100101111111" => data <= "000000";
				when "1100110000000" => data <= "000000";
				when "1100110000001" => data <= "000000";
				when "1100110000010" => data <= "000000";
				when "1100110000011" => data <= "000000";
				when "1100110000100" => data <= "000000";
				when "1100110000101" => data <= "000000";
				when "1100110000110" => data <= "000000";
				when "1100110000111" => data <= "000000";
				when "1100110001000" => data <= "000000";
				when "1100110001001" => data <= "000000";
				when "1100110001010" => data <= "000000";
				when "1100110001011" => data <= "000000";
				when "1100110001100" => data <= "000000";
				when "1100110001101" => data <= "000000";
				when "1100110001110" => data <= "000000";
				when "1100110001111" => data <= "000000";
				when "1100110010000" => data <= "000000";
				when "1100110010001" => data <= "000000";
				when "1100110010010" => data <= "000000";
				when "1100110010011" => data <= "000000";
				when "1100110010100" => data <= "000000";
				when "1100110010101" => data <= "000000";
				when "1100110010110" => data <= "000000";
				when "1100110010111" => data <= "000000";
				when "1100110011000" => data <= "000000";
				when "1100110011001" => data <= "000000";
				when "1100110011010" => data <= "000000";
				when "1100110011011" => data <= "000000";
				when "1100110011100" => data <= "000000";
				when "1100110011101" => data <= "000000";
				when "1100110011110" => data <= "000000";
				when "1100110011111" => data <= "000000";
				when "1100110100000" => data <= "000000";
				when "1100110100001" => data <= "000000";
				when "1100110100010" => data <= "000000";
				when "1100110100011" => data <= "000000";
				when "1100110100100" => data <= "000000";
				when "1100110100101" => data <= "000000";
				when "1100110100110" => data <= "000000";
				when "1100110100111" => data <= "000000";
				when "1100110101000" => data <= "000000";
				when "1100110101001" => data <= "000000";
				when "1100110101010" => data <= "000000";
				when "1100110101011" => data <= "000000";
				when "1100110101100" => data <= "000000";
				when "1100110101101" => data <= "000000";
				when "1100110101110" => data <= "000000";
				when "1100110101111" => data <= "010011";
				when "1100110110000" => data <= "010011";
				when "1100110110001" => data <= "010011";
				when "1100110110010" => data <= "010011";
				when "1100110110011" => data <= "010011";
				when "1100110110100" => data <= "000000";
				when "1100110110101" => data <= "000000";
				when "1100110110110" => data <= "000000";
				when "1100110110111" => data <= "000000";
				when "1100110111000" => data <= "000000";
				when "1100110111001" => data <= "000000";
				when "1100110111010" => data <= "000000";
				when "1100110111011" => data <= "000000";
				when "1100110111100" => data <= "000000";
				when "1100110111101" => data <= "000000";
				when "1100110111110" => data <= "000000";
				when "1100110111111" => data <= "000000";
				when "1100111000000" => data <= "000000";
				when "1100111000001" => data <= "000000";
				when "1100111000010" => data <= "000000";
				when "1100111000011" => data <= "000000";
				when "1100111000100" => data <= "000000";
				when "1100111000101" => data <= "000000";
				when "1100111000110" => data <= "000000";
				when "1100111000111" => data <= "000000";
				when "1100111001000" => data <= "000000";
				when "1100111001001" => data <= "000000";
				when "1100111001010" => data <= "000000";
				when "1100111001011" => data <= "000000";
				when "1100111001100" => data <= "000000";
				when "1100111001101" => data <= "000000";
				when "1100111001110" => data <= "000000";
				when "1100111001111" => data <= "000000";
				when "1100111010000" => data <= "000000";
				when "1100111010001" => data <= "010011";
				when "1100111010010" => data <= "000000";
				when "1100111010011" => data <= "000000";
				when "1100111010100" => data <= "000000";
				when "1100111010101" => data <= "000000";
				when "1100111010110" => data <= "000000";
				when "1100111010111" => data <= "000000";
				when "1100111011000" => data <= "000000";
				when "1100111011001" => data <= "000000";
				when "1100111011010" => data <= "000000";
				when "1100111011011" => data <= "000000";
				when "1100111011100" => data <= "000000";
				when "1100111011101" => data <= "000000";
				when "1100111011110" => data <= "000000";
				when "1100111011111" => data <= "000000";
				when "1100111100000" => data <= "000000";
				when "1100111100001" => data <= "000000";
				when "1100111100010" => data <= "000000";
				when "1100111100011" => data <= "000000";
				when "1100111100100" => data <= "000000";
				when "1100111100101" => data <= "000000";
				when "1100111100110" => data <= "000000";
				when "1100111100111" => data <= "000000";
				when "1100111101000" => data <= "000000";
				when "1100111101001" => data <= "000000";
				when "1100111101010" => data <= "000000";
				when "1100111101011" => data <= "000000";
				when "1100111101100" => data <= "000000";
				when "1100111101101" => data <= "000000";
				when "1100111101110" => data <= "000000";
				when "1100111101111" => data <= "000000";
				when "1100111110000" => data <= "000000";
				when "1100111110001" => data <= "000000";
				when "1100111110010" => data <= "000000";
				when "1100111110011" => data <= "000000";
				when "1100111110100" => data <= "000000";
				when "1100111110101" => data <= "000000";
				when "1100111110110" => data <= "000000";
				when "1100111110111" => data <= "000000";
				when "1100111111000" => data <= "000000";
				when "1100111111001" => data <= "000000";
				when "1100111111010" => data <= "000000";
				when "1100111111011" => data <= "000000";
				when "1100111111100" => data <= "000000";
				when "1100111111101" => data <= "000000";
				when "1100111111110" => data <= "000000";
				when "1100111111111" => data <= "000000";
				when "1101000000000" => data <= "000000";
				when "1101000000001" => data <= "000000";
				when "1101000000010" => data <= "000000";
				when "1101000000011" => data <= "000000";
				when "1101000000100" => data <= "000000";
				when "1101000000101" => data <= "000000";
				when "1101000000110" => data <= "000000";
				when "1101000000111" => data <= "000000";
				when "1101000001000" => data <= "000000";
				when "1101000001001" => data <= "000000";
				when "1101000001010" => data <= "000000";
				when "1101000001011" => data <= "000000";
				when "1101000001100" => data <= "000000";
				when "1101000001101" => data <= "000000";
				when "1101000001110" => data <= "000000";
				when "1101000001111" => data <= "000000";
				when "1101000010000" => data <= "000000";
				when "1101000010001" => data <= "000000";
				when "1101000010010" => data <= "000000";
				when "1101000010011" => data <= "000000";
				when "1101000010100" => data <= "000000";
				when "1101000010101" => data <= "000000";
				when "1101000010110" => data <= "000000";
				when "1101000010111" => data <= "000000";
				when "1101000011000" => data <= "000000";
				when "1101000011001" => data <= "000000";
				when "1101000011010" => data <= "000000";
				when "1101000011011" => data <= "000000";
				when "1101000011100" => data <= "000000";
				when "1101000011101" => data <= "000000";
				when "1101000011110" => data <= "000000";
				when "1101000011111" => data <= "000000";
				when "1101000100000" => data <= "000000";
				when "1101000100001" => data <= "000000";
				when "1101000100010" => data <= "000000";
				when "1101000100011" => data <= "000000";
				when "1101000100100" => data <= "000000";
				when "1101000100101" => data <= "000000";
				when "1101000100110" => data <= "000000";
				when "1101000100111" => data <= "000000";
				when "1101000101000" => data <= "000000";
				when "1101000101001" => data <= "000000";
				when "1101000101010" => data <= "000000";
				when "1101000101011" => data <= "000000";
				when "1101000101100" => data <= "000000";
				when "1101000101101" => data <= "000000";
				when "1101000101110" => data <= "000000";
				when "1101000101111" => data <= "010011";
				when "1101000110000" => data <= "000000";
				when "1101000110001" => data <= "000000";
				when "1101000110010" => data <= "000000";
				when "1101000110011" => data <= "010011";
				when "1101000110100" => data <= "010011";
				when "1101000110101" => data <= "000000";
				when "1101000110110" => data <= "000000";
				when "1101000110111" => data <= "000000";
				when "1101000111000" => data <= "000000";
				when "1101000111001" => data <= "000000";
				when "1101000111010" => data <= "000000";
				when "1101000111011" => data <= "000000";
				when "1101000111100" => data <= "000000";
				when "1101000111101" => data <= "000000";
				when "1101000111110" => data <= "000000";
				when "1101000111111" => data <= "000000";
				when "1101001000000" => data <= "000000";
				when "1101001000001" => data <= "000000";
				when "1101001000010" => data <= "000000";
				when "1101001000011" => data <= "000000";
				when "1101001000100" => data <= "000000";
				when "1101001000101" => data <= "000000";
				when "1101001000110" => data <= "000000";
				when "1101001000111" => data <= "000000";
				when "1101001001000" => data <= "000000";
				when "1101001001001" => data <= "000000";
				when "1101001001010" => data <= "000000";
				when "1101001001011" => data <= "000000";
				when "1101001001100" => data <= "000000";
				when "1101001001101" => data <= "000000";
				when "1101001001110" => data <= "000000";
				when "1101001001111" => data <= "000000";
				when "1101001010000" => data <= "000000";
				when "1101001010001" => data <= "010011";
				when "1101001010010" => data <= "000000";
				when "1101001010011" => data <= "000000";
				when "1101001010100" => data <= "000000";
				when "1101001010101" => data <= "000000";
				when "1101001010110" => data <= "000000";
				when "1101001010111" => data <= "000000";
				when "1101001011000" => data <= "000000";
				when "1101001011001" => data <= "000000";
				when "1101001011010" => data <= "000000";
				when "1101001011011" => data <= "000000";
				when "1101001011100" => data <= "000000";
				when "1101001011101" => data <= "000000";
				when "1101001011110" => data <= "000000";
				when "1101001011111" => data <= "000000";
				when "1101001100000" => data <= "000000";
				when "1101001100001" => data <= "000000";
				when "1101001100010" => data <= "000000";
				when "1101001100011" => data <= "000000";
				when "1101001100100" => data <= "000000";
				when "1101001100101" => data <= "000000";
				when "1101001100110" => data <= "000000";
				when "1101001100111" => data <= "000000";
				when "1101001101000" => data <= "000000";
				when "1101001101001" => data <= "000000";
				when "1101001101010" => data <= "000000";
				when "1101001101011" => data <= "000000";
				when "1101001101100" => data <= "000000";
				when "1101001101101" => data <= "000000";
				when "1101001101110" => data <= "000000";
				when "1101001101111" => data <= "000000";
				when "1101001110000" => data <= "000000";
				when "1101001110001" => data <= "000000";
				when "1101001110010" => data <= "000000";
				when "1101001110011" => data <= "000000";
				when "1101001110100" => data <= "000000";
				when "1101001110101" => data <= "000000";
				when "1101001110110" => data <= "000000";
				when "1101001110111" => data <= "000000";
				when "1101001111000" => data <= "000000";
				when "1101001111001" => data <= "000000";
				when "1101001111010" => data <= "000000";
				when "1101001111011" => data <= "000000";
				when "1101001111100" => data <= "000000";
				when "1101001111101" => data <= "000000";
				when "1101001111110" => data <= "000000";
				when "1101001111111" => data <= "000000";
				when "1101010000000" => data <= "000000";
				when "1101010000001" => data <= "000000";
				when "1101010000010" => data <= "000000";
				when "1101010000011" => data <= "000000";
				when "1101010000100" => data <= "000000";
				when "1101010000101" => data <= "000000";
				when "1101010000110" => data <= "000000";
				when "1101010000111" => data <= "000000";
				when "1101010001000" => data <= "000000";
				when "1101010001001" => data <= "000000";
				when "1101010001010" => data <= "000000";
				when "1101010001011" => data <= "000000";
				when "1101010001100" => data <= "000000";
				when "1101010001101" => data <= "000000";
				when "1101010001110" => data <= "000000";
				when "1101010001111" => data <= "000000";
				when "1101010010000" => data <= "000000";
				when "1101010010001" => data <= "000000";
				when "1101010010010" => data <= "000000";
				when "1101010010011" => data <= "000000";
				when "1101010010100" => data <= "000000";
				when "1101010010101" => data <= "000000";
				when "1101010010110" => data <= "000000";
				when "1101010010111" => data <= "000000";
				when "1101010011000" => data <= "000000";
				when "1101010011001" => data <= "000000";
				when "1101010011010" => data <= "000000";
				when "1101010011011" => data <= "000000";
				when "1101010011100" => data <= "000000";
				when "1101010011101" => data <= "000000";
				when "1101010011110" => data <= "000000";
				when "1101010011111" => data <= "000000";
				when "1101010100000" => data <= "000000";
				when "1101010100001" => data <= "000000";
				when "1101010100010" => data <= "000000";
				when "1101010100011" => data <= "000000";
				when "1101010100100" => data <= "000000";
				when "1101010100101" => data <= "000000";
				when "1101010100110" => data <= "000000";
				when "1101010100111" => data <= "000000";
				when "1101010101000" => data <= "000000";
				when "1101010101001" => data <= "000000";
				when "1101010101010" => data <= "000000";
				when "1101010101011" => data <= "000000";
				when "1101010101100" => data <= "000000";
				when "1101010101101" => data <= "000000";
				when "1101010101110" => data <= "000000";
				when "1101010101111" => data <= "010011";
				when "1101010110000" => data <= "000000";
				when "1101010110001" => data <= "000000";
				when "1101010110010" => data <= "000000";
				when "1101010110011" => data <= "010011";
				when "1101010110100" => data <= "010011";
				when "1101010110101" => data <= "000000";
				when "1101010110110" => data <= "000000";
				when "1101010110111" => data <= "000000";
				when "1101010111000" => data <= "000000";
				when "1101010111001" => data <= "000000";
				when "1101010111010" => data <= "000000";
				when "1101010111011" => data <= "000000";
				when "1101010111100" => data <= "010011";
				when "1101010111101" => data <= "010011";
				when "1101010111110" => data <= "010011";
				when "1101010111111" => data <= "010011";
				when "1101011000000" => data <= "010011";
				when "1101011000001" => data <= "010011";
				when "1101011000010" => data <= "010011";
				when "1101011000011" => data <= "010011";
				when "1101011000100" => data <= "010011";
				when "1101011000101" => data <= "010011";
				when "1101011000110" => data <= "000000";
				when "1101011000111" => data <= "000000";
				when "1101011001000" => data <= "000000";
				when "1101011001001" => data <= "000000";
				when "1101011001010" => data <= "000000";
				when "1101011001011" => data <= "000000";
				when "1101011001100" => data <= "000000";
				when "1101011001101" => data <= "000000";
				when "1101011001110" => data <= "000000";
				when "1101011001111" => data <= "000000";
				when "1101011010000" => data <= "000000";
				when "1101011010001" => data <= "010011";
				when "1101011010010" => data <= "000000";
				when "1101011010011" => data <= "000000";
				when "1101011010100" => data <= "000000";
				when "1101011010101" => data <= "000000";
				when "1101011010110" => data <= "000000";
				when "1101011010111" => data <= "000000";
				when "1101011011000" => data <= "000000";
				when "1101011011001" => data <= "000000";
				when "1101011011010" => data <= "000000";
				when "1101011011011" => data <= "000000";
				when "1101011011100" => data <= "000000";
				when "1101011011101" => data <= "000000";
				when "1101011011110" => data <= "000000";
				when "1101011011111" => data <= "000000";
				when "1101011100000" => data <= "000000";
				when "1101011100001" => data <= "000000";
				when "1101011100010" => data <= "000000";
				when "1101011100011" => data <= "000000";
				when "1101011100100" => data <= "000000";
				when "1101011100101" => data <= "000000";
				when "1101011100110" => data <= "000000";
				when "1101011100111" => data <= "000000";
				when "1101011101000" => data <= "000000";
				when "1101011101001" => data <= "000000";
				when "1101011101010" => data <= "000000";
				when "1101011101011" => data <= "000000";
				when "1101011101100" => data <= "000000";
				when "1101011101101" => data <= "000000";
				when "1101011101110" => data <= "000000";
				when "1101011101111" => data <= "000000";
				when "1101011110000" => data <= "000000";
				when "1101011110001" => data <= "000000";
				when "1101011110010" => data <= "000000";
				when "1101011110011" => data <= "000000";
				when "1101011110100" => data <= "000000";
				when "1101011110101" => data <= "000000";
				when "1101011110110" => data <= "000000";
				when "1101011110111" => data <= "000000";
				when "1101011111000" => data <= "000000";
				when "1101011111001" => data <= "000000";
				when "1101011111010" => data <= "000000";
				when "1101011111011" => data <= "000000";
				when "1101011111100" => data <= "000000";
				when "1101011111101" => data <= "000000";
				when "1101011111110" => data <= "000000";
				when "1101011111111" => data <= "000000";
				when "1101100000000" => data <= "000000";
				when "1101100000001" => data <= "000000";
				when "1101100000010" => data <= "000000";
				when "1101100000011" => data <= "000000";
				when "1101100000100" => data <= "000000";
				when "1101100000101" => data <= "000000";
				when "1101100000110" => data <= "000000";
				when "1101100000111" => data <= "000000";
				when "1101100001000" => data <= "000000";
				when "1101100001001" => data <= "000000";
				when "1101100001010" => data <= "000000";
				when "1101100001011" => data <= "000000";
				when "1101100001100" => data <= "000000";
				when "1101100001101" => data <= "000000";
				when "1101100001110" => data <= "000000";
				when "1101100001111" => data <= "000000";
				when "1101100010000" => data <= "000000";
				when "1101100010001" => data <= "000000";
				when "1101100010010" => data <= "000000";
				when "1101100010011" => data <= "000000";
				when "1101100010100" => data <= "000000";
				when "1101100010101" => data <= "000000";
				when "1101100010110" => data <= "000000";
				when "1101100010111" => data <= "000000";
				when "1101100011000" => data <= "000000";
				when "1101100011001" => data <= "000000";
				when "1101100011010" => data <= "000000";
				when "1101100011011" => data <= "000000";
				when "1101100011100" => data <= "000000";
				when "1101100011101" => data <= "000000";
				when "1101100011110" => data <= "000000";
				when "1101100011111" => data <= "000000";
				when "1101100100000" => data <= "000000";
				when "1101100100001" => data <= "000000";
				when "1101100100010" => data <= "000000";
				when "1101100100011" => data <= "000000";
				when "1101100100100" => data <= "000000";
				when "1101100100101" => data <= "000000";
				when "1101100100110" => data <= "000000";
				when "1101100100111" => data <= "000000";
				when "1101100101000" => data <= "000000";
				when "1101100101001" => data <= "000000";
				when "1101100101010" => data <= "000000";
				when "1101100101011" => data <= "000000";
				when "1101100101100" => data <= "000000";
				when "1101100101101" => data <= "000000";
				when "1101100101110" => data <= "000000";
				when "1101100101111" => data <= "010011";
				when "1101100110000" => data <= "000000";
				when "1101100110001" => data <= "000000";
				when "1101100110010" => data <= "000000";
				when "1101100110011" => data <= "000000";
				when "1101100110100" => data <= "010011";
				when "1101100110101" => data <= "010011";
				when "1101100110110" => data <= "000000";
				when "1101100110111" => data <= "000000";
				when "1101100111000" => data <= "000000";
				when "1101100111001" => data <= "000000";
				when "1101100111010" => data <= "000000";
				when "1101100111011" => data <= "000000";
				when "1101100111100" => data <= "010011";
				when "1101100111101" => data <= "000000";
				when "1101100111110" => data <= "000000";
				when "1101100111111" => data <= "000000";
				when "1101101000000" => data <= "000000";
				when "1101101000001" => data <= "000000";
				when "1101101000010" => data <= "000000";
				when "1101101000011" => data <= "000000";
				when "1101101000100" => data <= "000000";
				when "1101101000101" => data <= "010011";
				when "1101101000110" => data <= "000000";
				when "1101101000111" => data <= "000000";
				when "1101101001000" => data <= "000000";
				when "1101101001001" => data <= "000000";
				when "1101101001010" => data <= "000000";
				when "1101101001011" => data <= "000000";
				when "1101101001100" => data <= "000000";
				when "1101101001101" => data <= "000000";
				when "1101101001110" => data <= "000000";
				when "1101101001111" => data <= "000000";
				when "1101101010000" => data <= "000000";
				when "1101101010001" => data <= "010011";
				when "1101101010010" => data <= "000000";
				when "1101101010011" => data <= "000000";
				when "1101101010100" => data <= "000000";
				when "1101101010101" => data <= "000000";
				when "1101101010110" => data <= "000000";
				when "1101101010111" => data <= "000000";
				when "1101101011000" => data <= "000000";
				when "1101101011001" => data <= "000000";
				when "1101101011010" => data <= "000000";
				when "1101101011011" => data <= "000000";
				when "1101101011100" => data <= "000000";
				when "1101101011101" => data <= "000000";
				when "1101101011110" => data <= "000000";
				when "1101101011111" => data <= "000000";
				when "1101101100000" => data <= "000000";
				when "1101101100001" => data <= "000000";
				when "1101101100010" => data <= "000000";
				when "1101101100011" => data <= "000000";
				when "1101101100100" => data <= "000000";
				when "1101101100101" => data <= "000000";
				when "1101101100110" => data <= "000000";
				when "1101101100111" => data <= "000000";
				when "1101101101000" => data <= "000000";
				when "1101101101001" => data <= "000000";
				when "1101101101010" => data <= "000000";
				when "1101101101011" => data <= "000000";
				when "1101101101100" => data <= "000000";
				when "1101101101101" => data <= "000000";
				when "1101101101110" => data <= "000000";
				when "1101101101111" => data <= "000000";
				when "1101101110000" => data <= "000000";
				when "1101101110001" => data <= "000000";
				when "1101101110010" => data <= "000000";
				when "1101101110011" => data <= "000000";
				when "1101101110100" => data <= "000000";
				when "1101101110101" => data <= "000000";
				when "1101101110110" => data <= "000000";
				when "1101101110111" => data <= "000000";
				when "1101101111000" => data <= "000000";
				when "1101101111001" => data <= "000000";
				when "1101101111010" => data <= "000000";
				when "1101101111011" => data <= "000000";
				when "1101101111100" => data <= "000000";
				when "1101101111101" => data <= "000000";
				when "1101101111110" => data <= "000000";
				when "1101101111111" => data <= "000000";
				when "1101110000000" => data <= "000000";
				when "1101110000001" => data <= "000000";
				when "1101110000010" => data <= "000000";
				when "1101110000011" => data <= "000000";
				when "1101110000100" => data <= "000000";
				when "1101110000101" => data <= "000000";
				when "1101110000110" => data <= "000000";
				when "1101110000111" => data <= "000000";
				when "1101110001000" => data <= "000000";
				when "1101110001001" => data <= "000000";
				when "1101110001010" => data <= "000000";
				when "1101110001011" => data <= "000000";
				when "1101110001100" => data <= "000000";
				when "1101110001101" => data <= "000000";
				when "1101110001110" => data <= "000000";
				when "1101110001111" => data <= "000000";
				when "1101110010000" => data <= "000000";
				when "1101110010001" => data <= "000000";
				when "1101110010010" => data <= "000000";
				when "1101110010011" => data <= "000000";
				when "1101110010100" => data <= "000000";
				when "1101110010101" => data <= "000000";
				when "1101110010110" => data <= "000000";
				when "1101110010111" => data <= "000000";
				when "1101110011000" => data <= "000000";
				when "1101110011001" => data <= "000000";
				when "1101110011010" => data <= "000000";
				when "1101110011011" => data <= "000000";
				when "1101110011100" => data <= "000000";
				when "1101110011101" => data <= "000000";
				when "1101110011110" => data <= "000000";
				when "1101110011111" => data <= "000000";
				when "1101110100000" => data <= "000000";
				when "1101110100001" => data <= "000000";
				when "1101110100010" => data <= "000000";
				when "1101110100011" => data <= "000000";
				when "1101110100100" => data <= "000000";
				when "1101110100101" => data <= "000000";
				when "1101110100110" => data <= "000000";
				when "1101110100111" => data <= "000000";
				when "1101110101000" => data <= "000000";
				when "1101110101001" => data <= "000000";
				when "1101110101010" => data <= "000000";
				when "1101110101011" => data <= "000000";
				when "1101110101100" => data <= "000000";
				when "1101110101101" => data <= "000000";
				when "1101110101110" => data <= "000000";
				when "1101110101111" => data <= "010011";
				when "1101110110000" => data <= "000000";
				when "1101110110001" => data <= "000000";
				when "1101110110010" => data <= "000000";
				when "1101110110011" => data <= "000000";
				when "1101110110100" => data <= "010011";
				when "1101110110101" => data <= "010011";
				when "1101110110110" => data <= "000000";
				when "1101110110111" => data <= "000000";
				when "1101110111000" => data <= "000000";
				when "1101110111001" => data <= "000000";
				when "1101110111010" => data <= "000000";
				when "1101110111011" => data <= "000000";
				when "1101110111100" => data <= "010011";
				when "1101110111101" => data <= "010011";
				when "1101110111110" => data <= "010011";
				when "1101110111111" => data <= "010011";
				when "1101111000000" => data <= "010011";
				when "1101111000001" => data <= "010011";
				when "1101111000010" => data <= "010011";
				when "1101111000011" => data <= "010011";
				when "1101111000100" => data <= "010011";
				when "1101111000101" => data <= "010011";
				when "1101111000110" => data <= "000000";
				when "1101111000111" => data <= "000000";
				when "1101111001000" => data <= "000000";
				when "1101111001001" => data <= "000000";
				when "1101111001010" => data <= "000000";
				when "1101111001011" => data <= "000000";
				when "1101111001100" => data <= "000000";
				when "1101111001101" => data <= "000000";
				when "1101111001110" => data <= "000000";
				when "1101111001111" => data <= "000000";
				when "1101111010000" => data <= "000000";
				when "1101111010001" => data <= "010011";
				when "1101111010010" => data <= "000000";
				when "1101111010011" => data <= "000000";
				when "1101111010100" => data <= "000000";
				when "1101111010101" => data <= "000000";
				when "1101111010110" => data <= "000000";
				when "1101111010111" => data <= "000000";
				when "1101111011000" => data <= "000000";
				when "1101111011001" => data <= "000000";
				when "1101111011010" => data <= "000000";
				when "1101111011011" => data <= "000000";
				when "1101111011100" => data <= "000000";
				when "1101111011101" => data <= "000000";
				when "1101111011110" => data <= "000000";
				when "1101111011111" => data <= "000000";
				when "1101111100000" => data <= "000000";
				when "1101111100001" => data <= "000000";
				when "1101111100010" => data <= "000000";
				when "1101111100011" => data <= "000000";
				when "1101111100100" => data <= "000000";
				when "1101111100101" => data <= "000000";
				when "1101111100110" => data <= "000000";
				when "1101111100111" => data <= "000000";
				when "1101111101000" => data <= "000000";
				when "1101111101001" => data <= "000000";
				when "1101111101010" => data <= "000000";
				when "1101111101011" => data <= "000000";
				when "1101111101100" => data <= "000000";
				when "1101111101101" => data <= "000000";
				when "1101111101110" => data <= "000000";
				when "1101111101111" => data <= "000000";
				when "1101111110000" => data <= "000000";
				when "1101111110001" => data <= "000000";
				when "1101111110010" => data <= "000000";
				when "1101111110011" => data <= "000000";
				when "1101111110100" => data <= "000000";
				when "1101111110101" => data <= "000000";
				when "1101111110110" => data <= "000000";
				when "1101111110111" => data <= "000000";
				when "1101111111000" => data <= "000000";
				when "1101111111001" => data <= "000000";
				when "1101111111010" => data <= "000000";
				when "1101111111011" => data <= "000000";
				when "1101111111100" => data <= "000000";
				when "1101111111101" => data <= "000000";
				when "1101111111110" => data <= "000000";
				when "1101111111111" => data <= "000000";
				when "1110000000000" => data <= "000000";
				when "1110000000001" => data <= "000000";
				when "1110000000010" => data <= "000000";
				when "1110000000011" => data <= "000000";
				when "1110000000100" => data <= "000000";
				when "1110000000101" => data <= "000000";
				when "1110000000110" => data <= "000000";
				when "1110000000111" => data <= "000000";
				when "1110000001000" => data <= "000000";
				when "1110000001001" => data <= "000000";
				when "1110000001010" => data <= "000000";
				when "1110000001011" => data <= "000000";
				when "1110000001100" => data <= "000000";
				when "1110000001101" => data <= "000000";
				when "1110000001110" => data <= "000000";
				when "1110000001111" => data <= "000000";
				when "1110000010000" => data <= "000000";
				when "1110000010001" => data <= "000000";
				when "1110000010010" => data <= "000000";
				when "1110000010011" => data <= "000000";
				when "1110000010100" => data <= "000000";
				when "1110000010101" => data <= "000000";
				when "1110000010110" => data <= "000000";
				when "1110000010111" => data <= "000000";
				when "1110000011000" => data <= "000000";
				when "1110000011001" => data <= "000000";
				when "1110000011010" => data <= "000000";
				when "1110000011011" => data <= "000000";
				when "1110000011100" => data <= "000000";
				when "1110000011101" => data <= "000000";
				when "1110000011110" => data <= "000000";
				when "1110000011111" => data <= "000000";
				when "1110000100000" => data <= "000000";
				when "1110000100001" => data <= "000000";
				when "1110000100010" => data <= "000000";
				when "1110000100011" => data <= "000000";
				when "1110000100100" => data <= "000000";
				when "1110000100101" => data <= "000000";
				when "1110000100110" => data <= "000000";
				when "1110000100111" => data <= "000000";
				when "1110000101000" => data <= "000000";
				when "1110000101001" => data <= "000000";
				when "1110000101010" => data <= "000000";
				when "1110000101011" => data <= "000000";
				when "1110000101100" => data <= "000000";
				when "1110000101101" => data <= "000000";
				when "1110000101110" => data <= "000000";
				when "1110000101111" => data <= "010011";
				when "1110000110000" => data <= "000000";
				when "1110000110001" => data <= "000000";
				when "1110000110010" => data <= "000000";
				when "1110000110011" => data <= "000000";
				when "1110000110100" => data <= "010011";
				when "1110000110101" => data <= "000000";
				when "1110000110110" => data <= "000000";
				when "1110000110111" => data <= "000000";
				when "1110000111000" => data <= "000000";
				when "1110000111001" => data <= "000000";
				when "1110000111010" => data <= "000000";
				when "1110000111011" => data <= "000000";
				when "1110000111100" => data <= "010011";
				when "1110000111101" => data <= "000000";
				when "1110000111110" => data <= "000000";
				when "1110000111111" => data <= "000000";
				when "1110001000000" => data <= "000000";
				when "1110001000001" => data <= "000000";
				when "1110001000010" => data <= "000000";
				when "1110001000011" => data <= "000000";
				when "1110001000100" => data <= "000000";
				when "1110001000101" => data <= "010011";
				when "1110001000110" => data <= "000000";
				when "1110001000111" => data <= "000000";
				when "1110001001000" => data <= "000000";
				when "1110001001001" => data <= "000000";
				when "1110001001010" => data <= "000000";
				when "1110001001011" => data <= "000000";
				when "1110001001100" => data <= "000000";
				when "1110001001101" => data <= "000000";
				when "1110001001110" => data <= "000000";
				when "1110001001111" => data <= "000000";
				when "1110001010000" => data <= "000000";
				when "1110001010001" => data <= "010011";
				when "1110001010010" => data <= "000000";
				when "1110001010011" => data <= "000000";
				when "1110001010100" => data <= "000000";
				when "1110001010101" => data <= "000000";
				when "1110001010110" => data <= "000000";
				when "1110001010111" => data <= "000000";
				when "1110001011000" => data <= "000000";
				when "1110001011001" => data <= "000000";
				when "1110001011010" => data <= "000000";
				when "1110001011011" => data <= "000000";
				when "1110001011100" => data <= "000000";
				when "1110001011101" => data <= "000000";
				when "1110001011110" => data <= "000000";
				when "1110001011111" => data <= "000000";
				when "1110001100000" => data <= "000000";
				when "1110001100001" => data <= "000000";
				when "1110001100010" => data <= "000000";
				when "1110001100011" => data <= "000000";
				when "1110001100100" => data <= "000000";
				when "1110001100101" => data <= "000000";
				when "1110001100110" => data <= "000000";
				when "1110001100111" => data <= "000000";
				when "1110001101000" => data <= "000000";
				when "1110001101001" => data <= "000000";
				when "1110001101010" => data <= "000000";
				when "1110001101011" => data <= "000000";
				when "1110001101100" => data <= "000000";
				when "1110001101101" => data <= "000000";
				when "1110001101110" => data <= "000000";
				when "1110001101111" => data <= "000000";
				when "1110001110000" => data <= "000000";
				when "1110001110001" => data <= "000000";
				when "1110001110010" => data <= "000000";
				when "1110001110011" => data <= "000000";
				when "1110001110100" => data <= "000000";
				when "1110001110101" => data <= "000000";
				when "1110001110110" => data <= "000000";
				when "1110001110111" => data <= "000000";
				when "1110001111000" => data <= "000000";
				when "1110001111001" => data <= "000000";
				when "1110001111010" => data <= "000000";
				when "1110001111011" => data <= "000000";
				when "1110001111100" => data <= "000000";
				when "1110001111101" => data <= "000000";
				when "1110001111110" => data <= "000000";
				when "1110001111111" => data <= "000000";
				when "1110010000000" => data <= "000000";
				when "1110010000001" => data <= "000000";
				when "1110010000010" => data <= "000000";
				when "1110010000011" => data <= "000000";
				when "1110010000100" => data <= "000000";
				when "1110010000101" => data <= "000000";
				when "1110010000110" => data <= "000000";
				when "1110010000111" => data <= "000000";
				when "1110010001000" => data <= "000000";
				when "1110010001001" => data <= "000000";
				when "1110010001010" => data <= "000000";
				when "1110010001011" => data <= "000000";
				when "1110010001100" => data <= "000000";
				when "1110010001101" => data <= "000000";
				when "1110010001110" => data <= "000000";
				when "1110010001111" => data <= "000000";
				when "1110010010000" => data <= "000000";
				when "1110010010001" => data <= "000000";
				when "1110010010010" => data <= "000000";
				when "1110010010011" => data <= "000000";
				when "1110010010100" => data <= "000000";
				when "1110010010101" => data <= "000000";
				when "1110010010110" => data <= "000000";
				when "1110010010111" => data <= "000000";
				when "1110010011000" => data <= "000000";
				when "1110010011001" => data <= "000000";
				when "1110010011010" => data <= "000000";
				when "1110010011011" => data <= "000000";
				when "1110010011100" => data <= "000000";
				when "1110010011101" => data <= "000000";
				when "1110010011110" => data <= "000000";
				when "1110010011111" => data <= "000000";
				when "1110010100000" => data <= "000000";
				when "1110010100001" => data <= "000000";
				when "1110010100010" => data <= "000000";
				when "1110010100011" => data <= "000000";
				when "1110010100100" => data <= "000000";
				when "1110010100101" => data <= "000000";
				when "1110010100110" => data <= "000000";
				when "1110010100111" => data <= "000000";
				when "1110010101000" => data <= "000000";
				when "1110010101001" => data <= "000000";
				when "1110010101010" => data <= "000000";
				when "1110010101011" => data <= "000000";
				when "1110010101100" => data <= "000000";
				when "1110010101101" => data <= "000000";
				when "1110010101110" => data <= "000000";
				when "1110010101111" => data <= "010011";
				when "1110010110000" => data <= "000000";
				when "1110010110001" => data <= "000000";
				when "1110010110010" => data <= "000000";
				when "1110010110011" => data <= "010011";
				when "1110010110100" => data <= "000000";
				when "1110010110101" => data <= "000000";
				when "1110010110110" => data <= "000000";
				when "1110010110111" => data <= "000000";
				when "1110010111000" => data <= "000000";
				when "1110010111001" => data <= "000000";
				when "1110010111010" => data <= "000000";
				when "1110010111011" => data <= "000000";
				when "1110010111100" => data <= "010011";
				when "1110010111101" => data <= "000000";
				when "1110010111110" => data <= "000000";
				when "1110010111111" => data <= "000000";
				when "1110011000000" => data <= "000000";
				when "1110011000001" => data <= "000000";
				when "1110011000010" => data <= "000000";
				when "1110011000011" => data <= "000000";
				when "1110011000100" => data <= "000000";
				when "1110011000101" => data <= "010011";
				when "1110011000110" => data <= "000000";
				when "1110011000111" => data <= "000000";
				when "1110011001000" => data <= "000000";
				when "1110011001001" => data <= "000000";
				when "1110011001010" => data <= "000000";
				when "1110011001011" => data <= "000000";
				when "1110011001100" => data <= "000000";
				when "1110011001101" => data <= "000000";
				when "1110011001110" => data <= "000000";
				when "1110011001111" => data <= "000000";
				when "1110011010000" => data <= "000000";
				when "1110011010001" => data <= "010011";
				when "1110011010010" => data <= "000000";
				when "1110011010011" => data <= "000000";
				when "1110011010100" => data <= "000000";
				when "1110011010101" => data <= "000000";
				when "1110011010110" => data <= "000000";
				when "1110011010111" => data <= "000000";
				when "1110011011000" => data <= "000000";
				when "1110011011001" => data <= "000000";
				when "1110011011010" => data <= "000000";
				when "1110011011011" => data <= "000000";
				when "1110011011100" => data <= "000000";
				when "1110011011101" => data <= "000000";
				when "1110011011110" => data <= "000000";
				when "1110011011111" => data <= "000000";
				when "1110011100000" => data <= "000000";
				when "1110011100001" => data <= "000000";
				when "1110011100010" => data <= "000000";
				when "1110011100011" => data <= "000000";
				when "1110011100100" => data <= "000000";
				when "1110011100101" => data <= "000000";
				when "1110011100110" => data <= "000000";
				when "1110011100111" => data <= "000000";
				when "1110011101000" => data <= "000000";
				when "1110011101001" => data <= "000000";
				when "1110011101010" => data <= "000000";
				when "1110011101011" => data <= "000000";
				when "1110011101100" => data <= "000000";
				when "1110011101101" => data <= "000000";
				when "1110011101110" => data <= "000000";
				when "1110011101111" => data <= "000000";
				when "1110011110000" => data <= "000000";
				when "1110011110001" => data <= "000000";
				when "1110011110010" => data <= "000000";
				when "1110011110011" => data <= "000000";
				when "1110011110100" => data <= "000000";
				when "1110011110101" => data <= "000000";
				when "1110011110110" => data <= "000000";
				when "1110011110111" => data <= "000000";
				when "1110011111000" => data <= "000000";
				when "1110011111001" => data <= "000000";
				when "1110011111010" => data <= "000000";
				when "1110011111011" => data <= "000000";
				when "1110011111100" => data <= "000000";
				when "1110011111101" => data <= "000000";
				when "1110011111110" => data <= "000000";
				when "1110011111111" => data <= "000000";
				when "1110100000000" => data <= "000000";
				when "1110100000001" => data <= "000000";
				when "1110100000010" => data <= "000000";
				when "1110100000011" => data <= "000000";
				when "1110100000100" => data <= "000000";
				when "1110100000101" => data <= "000000";
				when "1110100000110" => data <= "000000";
				when "1110100000111" => data <= "000000";
				when "1110100001000" => data <= "000000";
				when "1110100001001" => data <= "000000";
				when "1110100001010" => data <= "000000";
				when "1110100001011" => data <= "000000";
				when "1110100001100" => data <= "000000";
				when "1110100001101" => data <= "000000";
				when "1110100001110" => data <= "000000";
				when "1110100001111" => data <= "000000";
				when "1110100010000" => data <= "000000";
				when "1110100010001" => data <= "000000";
				when "1110100010010" => data <= "000000";
				when "1110100010011" => data <= "000000";
				when "1110100010100" => data <= "000000";
				when "1110100010101" => data <= "000000";
				when "1110100010110" => data <= "000000";
				when "1110100010111" => data <= "000000";
				when "1110100011000" => data <= "000000";
				when "1110100011001" => data <= "000000";
				when "1110100011010" => data <= "000000";
				when "1110100011011" => data <= "000000";
				when "1110100011100" => data <= "000000";
				when "1110100011101" => data <= "000000";
				when "1110100011110" => data <= "000000";
				when "1110100011111" => data <= "000000";
				when "1110100100000" => data <= "000000";
				when "1110100100001" => data <= "000000";
				when "1110100100010" => data <= "000000";
				when "1110100100011" => data <= "000000";
				when "1110100100100" => data <= "000000";
				when "1110100100101" => data <= "000000";
				when "1110100100110" => data <= "000000";
				when "1110100100111" => data <= "000000";
				when "1110100101000" => data <= "000000";
				when "1110100101001" => data <= "000000";
				when "1110100101010" => data <= "000000";
				when "1110100101011" => data <= "000000";
				when "1110100101100" => data <= "000000";
				when "1110100101101" => data <= "000000";
				when "1110100101110" => data <= "000000";
				when "1110100101111" => data <= "010011";
				when "1110100110000" => data <= "000000";
				when "1110100110001" => data <= "000000";
				when "1110100110010" => data <= "000000";
				when "1110100110011" => data <= "000000";
				when "1110100110100" => data <= "000000";
				when "1110100110101" => data <= "000000";
				when "1110100110110" => data <= "000000";
				when "1110100110111" => data <= "000000";
				when "1110100111000" => data <= "000000";
				when "1110100111001" => data <= "000000";
				when "1110100111010" => data <= "000000";
				when "1110100111011" => data <= "000000";
				when "1110100111100" => data <= "010011";
				when "1110100111101" => data <= "000000";
				when "1110100111110" => data <= "000000";
				when "1110100111111" => data <= "000000";
				when "1110101000000" => data <= "000000";
				when "1110101000001" => data <= "000000";
				when "1110101000010" => data <= "000000";
				when "1110101000011" => data <= "000000";
				when "1110101000100" => data <= "000000";
				when "1110101000101" => data <= "010011";
				when "1110101000110" => data <= "000000";
				when "1110101000111" => data <= "000000";
				when "1110101001000" => data <= "000000";
				when "1110101001001" => data <= "000000";
				when "1110101001010" => data <= "000000";
				when "1110101001011" => data <= "000000";
				when "1110101001100" => data <= "000000";
				when "1110101001101" => data <= "000000";
				when "1110101001110" => data <= "000000";
				when "1110101001111" => data <= "000000";
				when "1110101010000" => data <= "000000";
				when "1110101010001" => data <= "010011";
				when "1110101010010" => data <= "000000";
				when "1110101010011" => data <= "000000";
				when "1110101010100" => data <= "000000";
				when "1110101010101" => data <= "000000";
				when "1110101010110" => data <= "000000";
				when "1110101010111" => data <= "000000";
				when "1110101011000" => data <= "000000";
				when "1110101011001" => data <= "000000";
				when "1110101011010" => data <= "000000";
				when "1110101011011" => data <= "000000";
				when "1110101011100" => data <= "000000";
				when "1110101011101" => data <= "000000";
				when "1110101011110" => data <= "000000";
				when "1110101011111" => data <= "000000";
				when "1110101100000" => data <= "000000";
				when "1110101100001" => data <= "000000";
				when "1110101100010" => data <= "000000";
				when "1110101100011" => data <= "000000";
				when "1110101100100" => data <= "000000";
				when "1110101100101" => data <= "000000";
				when "1110101100110" => data <= "000000";
				when "1110101100111" => data <= "000000";
				when "1110101101000" => data <= "000000";
				when "1110101101001" => data <= "000000";
				when "1110101101010" => data <= "000000";
				when "1110101101011" => data <= "000000";
				when "1110101101100" => data <= "000000";
				when "1110101101101" => data <= "000000";
				when "1110101101110" => data <= "000000";
				when "1110101101111" => data <= "000000";
				when "1110101110000" => data <= "000000";
				when "1110101110001" => data <= "000000";
				when "1110101110010" => data <= "000000";
				when "1110101110011" => data <= "000000";
				when "1110101110100" => data <= "000000";
				when "1110101110101" => data <= "000000";
				when "1110101110110" => data <= "000000";
				when "1110101110111" => data <= "000000";
				when "1110101111000" => data <= "000000";
				when "1110101111001" => data <= "000000";
				when "1110101111010" => data <= "000000";
				when "1110101111011" => data <= "000000";
				when "1110101111100" => data <= "000000";
				when "1110101111101" => data <= "000000";
				when "1110101111110" => data <= "000000";
				when "1110101111111" => data <= "000000";
				when "1110110000000" => data <= "000000";
				when "1110110000001" => data <= "000000";
				when "1110110000010" => data <= "000000";
				when "1110110000011" => data <= "000000";
				when "1110110000100" => data <= "000000";
				when "1110110000101" => data <= "000000";
				when "1110110000110" => data <= "000000";
				when "1110110000111" => data <= "000000";
				when "1110110001000" => data <= "000000";
				when "1110110001001" => data <= "000000";
				when "1110110001010" => data <= "000000";
				when "1110110001011" => data <= "000000";
				when "1110110001100" => data <= "000000";
				when "1110110001101" => data <= "000000";
				when "1110110001110" => data <= "000000";
				when "1110110001111" => data <= "000000";
				when "1110110010000" => data <= "000000";
				when "1110110010001" => data <= "000000";
				when "1110110010010" => data <= "000000";
				when "1110110010011" => data <= "000000";
				when "1110110010100" => data <= "000000";
				when "1110110010101" => data <= "000000";
				when "1110110010110" => data <= "000000";
				when "1110110010111" => data <= "000000";
				when "1110110011000" => data <= "000000";
				when "1110110011001" => data <= "000000";
				when "1110110011010" => data <= "000000";
				when "1110110011011" => data <= "000000";
				when "1110110011100" => data <= "000000";
				when "1110110011101" => data <= "000000";
				when "1110110011110" => data <= "000000";
				when "1110110011111" => data <= "000000";
				when "1110110100000" => data <= "000000";
				when "1110110100001" => data <= "000000";
				when "1110110100010" => data <= "000000";
				when "1110110100011" => data <= "000000";
				when "1110110100100" => data <= "000000";
				when "1110110100101" => data <= "000000";
				when "1110110100110" => data <= "000000";
				when "1110110100111" => data <= "000000";
				when "1110110101000" => data <= "000000";
				when "1110110101001" => data <= "000000";
				when "1110110101010" => data <= "000000";
				when "1110110101011" => data <= "000000";
				when "1110110101100" => data <= "000000";
				when "1110110101101" => data <= "000000";
				when "1110110101110" => data <= "000000";
				when "1110110101111" => data <= "010011";
				when "1110110110000" => data <= "000000";
				when "1110110110001" => data <= "000000";
				when "1110110110010" => data <= "000000";
				when "1110110110011" => data <= "000000";
				when "1110110110100" => data <= "000000";
				when "1110110110101" => data <= "000000";
				when "1110110110110" => data <= "000000";
				when "1110110110111" => data <= "000000";
				when "1110110111000" => data <= "000000";
				when "1110110111001" => data <= "000000";
				when "1110110111010" => data <= "000000";
				when "1110110111011" => data <= "000000";
				when "1110110111100" => data <= "010011";
				when "1110110111101" => data <= "000000";
				when "1110110111110" => data <= "000000";
				when "1110110111111" => data <= "000000";
				when "1110111000000" => data <= "000000";
				when "1110111000001" => data <= "000000";
				when "1110111000010" => data <= "000000";
				when "1110111000011" => data <= "000000";
				when "1110111000100" => data <= "000000";
				when "1110111000101" => data <= "010011";
				when "1110111000110" => data <= "000000";
				when "1110111000111" => data <= "000000";
				when "1110111001000" => data <= "000000";
				when "1110111001001" => data <= "000000";
				when "1110111001010" => data <= "000000";
				when "1110111001011" => data <= "000000";
				when "1110111001100" => data <= "010011";
				when "1110111001101" => data <= "010011";
				when "1110111001110" => data <= "010011";
				when "1110111001111" => data <= "010011";
				when "1110111010000" => data <= "010011";
				when "1110111010001" => data <= "010011";
				when "1110111010010" => data <= "000000";
				when "1110111010011" => data <= "000000";
				when "1110111010100" => data <= "000000";
				when "1110111010101" => data <= "000000";
				when "1110111010110" => data <= "000000";
				when "1110111010111" => data <= "000000";
				when "1110111011000" => data <= "000000";
				when "1110111011001" => data <= "000000";
				when "1110111011010" => data <= "000000";
				when "1110111011011" => data <= "000000";
				when "1110111011100" => data <= "000000";
				when "1110111011101" => data <= "000000";
				when "1110111011110" => data <= "000000";
				when "1110111011111" => data <= "000000";
				when "1110111100000" => data <= "000000";
				when "1110111100001" => data <= "000000";
				when "1110111100010" => data <= "000000";
				when "1110111100011" => data <= "000000";
				when "1110111100100" => data <= "000000";
				when "1110111100101" => data <= "000000";
				when "1110111100110" => data <= "000000";
				when "1110111100111" => data <= "000000";
				when "1110111101000" => data <= "000000";
				when "1110111101001" => data <= "000000";
				when "1110111101010" => data <= "000000";
				when "1110111101011" => data <= "000000";
				when "1110111101100" => data <= "000000";
				when "1110111101101" => data <= "000000";
				when "1110111101110" => data <= "000000";
				when "1110111101111" => data <= "000000";
				when "1110111110000" => data <= "000000";
				when "1110111110001" => data <= "000000";
				when "1110111110010" => data <= "000000";
				when "1110111110011" => data <= "000000";
				when "1110111110100" => data <= "000000";
				when "1110111110101" => data <= "000000";
				when "1110111110110" => data <= "000000";
				when "1110111110111" => data <= "000000";
				when "1110111111000" => data <= "000000";
				when "1110111111001" => data <= "000000";
				when "1110111111010" => data <= "000000";
				when "1110111111011" => data <= "000000";
				when "1110111111100" => data <= "000000";
				when "1110111111101" => data <= "000000";
				when "1110111111110" => data <= "000000";
				when "1110111111111" => data <= "000000";
				when "1111000000000" => data <= "000000";
				when "1111000000001" => data <= "000000";
				when "1111000000010" => data <= "000000";
				when "1111000000011" => data <= "000000";
				when "1111000000100" => data <= "000000";
				when "1111000000101" => data <= "000000";
				when "1111000000110" => data <= "000000";
				when "1111000000111" => data <= "000000";
				when "1111000001000" => data <= "000000";
				when "1111000001001" => data <= "000000";
				when "1111000001010" => data <= "000000";
				when "1111000001011" => data <= "000000";
				when "1111000001100" => data <= "000000";
				when "1111000001101" => data <= "000000";
				when "1111000001110" => data <= "000000";
				when "1111000001111" => data <= "000000";
				when "1111000010000" => data <= "000000";
				when "1111000010001" => data <= "000000";
				when "1111000010010" => data <= "000000";
				when "1111000010011" => data <= "000000";
				when "1111000010100" => data <= "000000";
				when "1111000010101" => data <= "000000";
				when "1111000010110" => data <= "000000";
				when "1111000010111" => data <= "000000";
				when "1111000011000" => data <= "000000";
				when "1111000011001" => data <= "000000";
				when "1111000011010" => data <= "000000";
				when "1111000011011" => data <= "000000";
				when "1111000011100" => data <= "000000";
				when "1111000011101" => data <= "000000";
				when "1111000011110" => data <= "000000";
				when "1111000011111" => data <= "000000";
				when "1111000100000" => data <= "000000";
				when "1111000100001" => data <= "000000";
				when "1111000100010" => data <= "000000";
				when "1111000100011" => data <= "000000";
				when "1111000100100" => data <= "000000";
				when "1111000100101" => data <= "000000";
				when "1111000100110" => data <= "000000";
				when "1111000100111" => data <= "000000";
				when "1111000101000" => data <= "000000";
				when "1111000101001" => data <= "000000";
				when "1111000101010" => data <= "000000";
				when "1111000101011" => data <= "010011";
				when "1111000101100" => data <= "010011";
				when "1111000101101" => data <= "010011";
				when "1111000101110" => data <= "010011";
				when "1111000101111" => data <= "010011";
				when "1111000110000" => data <= "000000";
				when "1111000110001" => data <= "000000";
				when "1111000110010" => data <= "000000";
				when "1111000110011" => data <= "000000";
				when "1111000110100" => data <= "000000";
				when "1111000110101" => data <= "000000";
				when "1111000110110" => data <= "000000";
				when "1111000110111" => data <= "000000";
				when "1111000111000" => data <= "000000";
				when "1111000111001" => data <= "000000";
				when "1111000111010" => data <= "000000";
				when "1111000111011" => data <= "000000";
				when "1111000111100" => data <= "010011";
				when "1111000111101" => data <= "000000";
				when "1111000111110" => data <= "000000";
				when "1111000111111" => data <= "000000";
				when "1111001000000" => data <= "000000";
				when "1111001000001" => data <= "000000";
				when "1111001000010" => data <= "000000";
				when "1111001000011" => data <= "000000";
				when "1111001000100" => data <= "000000";
				when "1111001000101" => data <= "010011";
				when "1111001000110" => data <= "000000";
				when "1111001000111" => data <= "000000";
				when "1111001001000" => data <= "000000";
				when "1111001001001" => data <= "000000";
				when "1111001001010" => data <= "000000";
				when "1111001001011" => data <= "010011";
				when "1111001001100" => data <= "010011";
				when "1111001001101" => data <= "010011";
				when "1111001001110" => data <= "010011";
				when "1111001001111" => data <= "010011";
				when "1111001010000" => data <= "010011";
				when "1111001010001" => data <= "010011";
				when "1111001010010" => data <= "000000";
				when "1111001010011" => data <= "000000";
				when "1111001010100" => data <= "000000";
				when "1111001010101" => data <= "000000";
				when "1111001010110" => data <= "000000";
				when "1111001010111" => data <= "000000";
				when "1111001011000" => data <= "000000";
				when "1111001011001" => data <= "000000";
				when "1111001011010" => data <= "000000";
				when "1111001011011" => data <= "000000";
				when "1111001011100" => data <= "000000";
				when "1111001011101" => data <= "000000";
				when "1111001011110" => data <= "000000";
				when "1111001011111" => data <= "000000";
				when "1111001100000" => data <= "000000";
				when "1111001100001" => data <= "000000";
				when "1111001100010" => data <= "000000";
				when "1111001100011" => data <= "000000";
				when "1111001100100" => data <= "000000";
				when "1111001100101" => data <= "000000";
				when "1111001100110" => data <= "000000";
				when "1111001100111" => data <= "000000";
				when "1111001101000" => data <= "000000";
				when "1111001101001" => data <= "000000";
				when "1111001101010" => data <= "000000";
				when "1111001101011" => data <= "000000";
				when "1111001101100" => data <= "000000";
				when "1111001101101" => data <= "000000";
				when "1111001101110" => data <= "000000";
				when "1111001101111" => data <= "000000";
				when "1111001110000" => data <= "000000";
				when "1111001110001" => data <= "000000";
				when "1111001110010" => data <= "000000";
				when "1111001110011" => data <= "000000";
				when "1111001110100" => data <= "000000";
				when "1111001110101" => data <= "000000";
				when "1111001110110" => data <= "000000";
				when "1111001110111" => data <= "000000";
				when "1111001111000" => data <= "000000";
				when "1111001111001" => data <= "000000";
				when "1111001111010" => data <= "000000";
				when "1111001111011" => data <= "000000";
				when "1111001111100" => data <= "000000";
				when "1111001111101" => data <= "000000";
				when "1111001111110" => data <= "000000";
				when "1111001111111" => data <= "000000";
				when "1111010000000" => data <= "000000";
				when "1111010000001" => data <= "000000";
				when "1111010000010" => data <= "000000";
				when "1111010000011" => data <= "000000";
				when "1111010000100" => data <= "000000";
				when "1111010000101" => data <= "000000";
				when "1111010000110" => data <= "000000";
				when "1111010000111" => data <= "000000";
				when "1111010001000" => data <= "000000";
				when "1111010001001" => data <= "000000";
				when "1111010001010" => data <= "000000";
				when "1111010001011" => data <= "000000";
				when "1111010001100" => data <= "000000";
				when "1111010001101" => data <= "000000";
				when "1111010001110" => data <= "000000";
				when "1111010001111" => data <= "000000";
				when "1111010010000" => data <= "000000";
				when "1111010010001" => data <= "000000";
				when "1111010010010" => data <= "000000";
				when "1111010010011" => data <= "000000";
				when "1111010010100" => data <= "000000";
				when "1111010010101" => data <= "000000";
				when "1111010010110" => data <= "000000";
				when "1111010010111" => data <= "000000";
				when "1111010011000" => data <= "000000";
				when "1111010011001" => data <= "000000";
				when "1111010011010" => data <= "000000";
				when "1111010011011" => data <= "000000";
				when "1111010011100" => data <= "000000";
				when "1111010011101" => data <= "000000";
				when "1111010011110" => data <= "000000";
				when "1111010011111" => data <= "000000";
				when "1111010100000" => data <= "000000";
				when "1111010100001" => data <= "000000";
				when "1111010100010" => data <= "000000";
				when "1111010100011" => data <= "000000";
				when "1111010100100" => data <= "000000";
				when "1111010100101" => data <= "000000";
				when "1111010100110" => data <= "000000";
				when "1111010100111" => data <= "000000";
				when "1111010101000" => data <= "000000";
				when "1111010101001" => data <= "000000";
				when "1111010101010" => data <= "010011";
				when "1111010101011" => data <= "010011";
				when "1111010101100" => data <= "010011";
				when "1111010101101" => data <= "010011";
				when "1111010101110" => data <= "010011";
				when "1111010101111" => data <= "010011";
				when "1111010110000" => data <= "000000";
				when "1111010110001" => data <= "000000";
				when "1111010110010" => data <= "000000";
				when "1111010110011" => data <= "000000";
				when "1111010110100" => data <= "000000";
				when "1111010110101" => data <= "000000";
				when "1111010110110" => data <= "000000";
				when "1111010110111" => data <= "000000";
				when "1111010111000" => data <= "010011";
				when "1111010111001" => data <= "010011";
				when "1111010111010" => data <= "010011";
				when "1111010111011" => data <= "010011";
				when "1111010111100" => data <= "010011";
				when "1111010111101" => data <= "000000";
				when "1111010111110" => data <= "000000";
				when "1111010111111" => data <= "000000";
				when "1111011000000" => data <= "000000";
				when "1111011000001" => data <= "010011";
				when "1111011000010" => data <= "010011";
				when "1111011000011" => data <= "010011";
				when "1111011000100" => data <= "010011";
				when "1111011000101" => data <= "010011";
				when "1111011000110" => data <= "000000";
				when "1111011000111" => data <= "000000";
				when "1111011001000" => data <= "000000";
				when "1111011001001" => data <= "000000";
				when "1111011001010" => data <= "000000";
				when "1111011001011" => data <= "010011";
				when "1111011001100" => data <= "111111";
				when "1111011001101" => data <= "010011";
				when "1111011001110" => data <= "010011";
				when "1111011001111" => data <= "010011";
				when "1111011010000" => data <= "010011";
				when "1111011010001" => data <= "010011";
				when "1111011010010" => data <= "000000";
				when "1111011010011" => data <= "000000";
				when "1111011010100" => data <= "000000";
				when "1111011010101" => data <= "000000";
				when "1111011010110" => data <= "000000";
				when "1111011010111" => data <= "000000";
				when "1111011011000" => data <= "000000";
				when "1111011011001" => data <= "000000";
				when "1111011011010" => data <= "000000";
				when "1111011011011" => data <= "000000";
				when "1111011011100" => data <= "000000";
				when "1111011011101" => data <= "000000";
				when "1111011011110" => data <= "000000";
				when "1111011011111" => data <= "000000";
				when "1111011100000" => data <= "000000";
				when "1111011100001" => data <= "000000";
				when "1111011100010" => data <= "000000";
				when "1111011100011" => data <= "000000";
				when "1111011100100" => data <= "000000";
				when "1111011100101" => data <= "000000";
				when "1111011100110" => data <= "000000";
				when "1111011100111" => data <= "000000";
				when "1111011101000" => data <= "000000";
				when "1111011101001" => data <= "000000";
				when "1111011101010" => data <= "000000";
				when "1111011101011" => data <= "000000";
				when "1111011101100" => data <= "000000";
				when "1111011101101" => data <= "000000";
				when "1111011101110" => data <= "000000";
				when "1111011101111" => data <= "000000";
				when "1111011110000" => data <= "000000";
				when "1111011110001" => data <= "000000";
				when "1111011110010" => data <= "000000";
				when "1111011110011" => data <= "000000";
				when "1111011110100" => data <= "000000";
				when "1111011110101" => data <= "000000";
				when "1111011110110" => data <= "000000";
				when "1111011110111" => data <= "000000";
				when "1111011111000" => data <= "000000";
				when "1111011111001" => data <= "000000";
				when "1111011111010" => data <= "000000";
				when "1111011111011" => data <= "000000";
				when "1111011111100" => data <= "000000";
				when "1111011111101" => data <= "000000";
				when "1111011111110" => data <= "000000";
				when "1111011111111" => data <= "000000";
				when "1111100000000" => data <= "000000";
				when "1111100000001" => data <= "000000";
				when "1111100000010" => data <= "000000";
				when "1111100000011" => data <= "000000";
				when "1111100000100" => data <= "000000";
				when "1111100000101" => data <= "000000";
				when "1111100000110" => data <= "000000";
				when "1111100000111" => data <= "000000";
				when "1111100001000" => data <= "000000";
				when "1111100001001" => data <= "000000";
				when "1111100001010" => data <= "000000";
				when "1111100001011" => data <= "000000";
				when "1111100001100" => data <= "000000";
				when "1111100001101" => data <= "000000";
				when "1111100001110" => data <= "000000";
				when "1111100001111" => data <= "000000";
				when "1111100010000" => data <= "000000";
				when "1111100010001" => data <= "000000";
				when "1111100010010" => data <= "000000";
				when "1111100010011" => data <= "000000";
				when "1111100010100" => data <= "000000";
				when "1111100010101" => data <= "000000";
				when "1111100010110" => data <= "000000";
				when "1111100010111" => data <= "000000";
				when "1111100011000" => data <= "000000";
				when "1111100011001" => data <= "000000";
				when "1111100011010" => data <= "000000";
				when "1111100011011" => data <= "000000";
				when "1111100011100" => data <= "000000";
				when "1111100011101" => data <= "000000";
				when "1111100011110" => data <= "000000";
				when "1111100011111" => data <= "000000";
				when "1111100100000" => data <= "000000";
				when "1111100100001" => data <= "000000";
				when "1111100100010" => data <= "000000";
				when "1111100100011" => data <= "000000";
				when "1111100100100" => data <= "000000";
				when "1111100100101" => data <= "000000";
				when "1111100100110" => data <= "000000";
				when "1111100100111" => data <= "000000";
				when "1111100101000" => data <= "000000";
				when "1111100101001" => data <= "000000";
				when "1111100101010" => data <= "010011";
				when "1111100101011" => data <= "111111";
				when "1111100101100" => data <= "010011";
				when "1111100101101" => data <= "010011";
				when "1111100101110" => data <= "010011";
				when "1111100101111" => data <= "010011";
				when "1111100110000" => data <= "000000";
				when "1111100110001" => data <= "000000";
				when "1111100110010" => data <= "000000";
				when "1111100110011" => data <= "000000";
				when "1111100110100" => data <= "000000";
				when "1111100110101" => data <= "000000";
				when "1111100110110" => data <= "000000";
				when "1111100110111" => data <= "010011";
				when "1111100111000" => data <= "010011";
				when "1111100111001" => data <= "010011";
				when "1111100111010" => data <= "010011";
				when "1111100111011" => data <= "010011";
				when "1111100111100" => data <= "010011";
				when "1111100111101" => data <= "000000";
				when "1111100111110" => data <= "000000";
				when "1111100111111" => data <= "000000";
				when "1111101000000" => data <= "010011";
				when "1111101000001" => data <= "010011";
				when "1111101000010" => data <= "010011";
				when "1111101000011" => data <= "010011";
				when "1111101000100" => data <= "010011";
				when "1111101000101" => data <= "010011";
				when "1111101000110" => data <= "000000";
				when "1111101000111" => data <= "000000";
				when "1111101001000" => data <= "000000";
				when "1111101001001" => data <= "000000";
				when "1111101001010" => data <= "000000";
				when "1111101001011" => data <= "010011";
				when "1111101001100" => data <= "010011";
				when "1111101001101" => data <= "010011";
				when "1111101001110" => data <= "010011";
				when "1111101001111" => data <= "010011";
				when "1111101010000" => data <= "010011";
				when "1111101010001" => data <= "010011";
				when "1111101010010" => data <= "000000";
				when "1111101010011" => data <= "000000";
				when "1111101010100" => data <= "000000";
				when "1111101010101" => data <= "000000";
				when "1111101010110" => data <= "000000";
				when "1111101010111" => data <= "000000";
				when "1111101011000" => data <= "000000";
				when "1111101011001" => data <= "000000";
				when "1111101011010" => data <= "000000";
				when "1111101011011" => data <= "000000";
				when "1111101011100" => data <= "000000";
				when "1111101011101" => data <= "000000";
				when "1111101011110" => data <= "000000";
				when "1111101011111" => data <= "000000";
				when "1111101100000" => data <= "000000";
				when "1111101100001" => data <= "000000";
				when "1111101100010" => data <= "000000";
				when "1111101100011" => data <= "000000";
				when "1111101100100" => data <= "000000";
				when "1111101100101" => data <= "000000";
				when "1111101100110" => data <= "000000";
				when "1111101100111" => data <= "000000";
				when "1111101101000" => data <= "000000";
				when "1111101101001" => data <= "000000";
				when "1111101101010" => data <= "000000";
				when "1111101101011" => data <= "000000";
				when "1111101101100" => data <= "000000";
				when "1111101101101" => data <= "000000";
				when "1111101101110" => data <= "000000";
				when "1111101101111" => data <= "000000";
				when "1111101110000" => data <= "000000";
				when "1111101110001" => data <= "000000";
				when "1111101110010" => data <= "000000";
				when "1111101110011" => data <= "000000";
				when "1111101110100" => data <= "000000";
				when "1111101110101" => data <= "000000";
				when "1111101110110" => data <= "000000";
				when "1111101110111" => data <= "000000";
				when "1111101111000" => data <= "000000";
				when "1111101111001" => data <= "000000";
				when "1111101111010" => data <= "000000";
				when "1111101111011" => data <= "000000";
				when "1111101111100" => data <= "000000";
				when "1111101111101" => data <= "000000";
				when "1111101111110" => data <= "000000";
				when "1111101111111" => data <= "000000";
				when "1111110000000" => data <= "000000";
				when "1111110000001" => data <= "000000";
				when "1111110000010" => data <= "000000";
				when "1111110000011" => data <= "000000";
				when "1111110000100" => data <= "000000";
				when "1111110000101" => data <= "000000";
				when "1111110000110" => data <= "000000";
				when "1111110000111" => data <= "000000";
				when "1111110001000" => data <= "000000";
				when "1111110001001" => data <= "000000";
				when "1111110001010" => data <= "000000";
				when "1111110001011" => data <= "000000";
				when "1111110001100" => data <= "000000";
				when "1111110001101" => data <= "000000";
				when "1111110001110" => data <= "000000";
				when "1111110001111" => data <= "000000";
				when "1111110010000" => data <= "000000";
				when "1111110010001" => data <= "000000";
				when "1111110010010" => data <= "000000";
				when "1111110010011" => data <= "000000";
				when "1111110010100" => data <= "000000";
				when "1111110010101" => data <= "000000";
				when "1111110010110" => data <= "000000";
				when "1111110010111" => data <= "000000";
				when "1111110011000" => data <= "000000";
				when "1111110011001" => data <= "000000";
				when "1111110011010" => data <= "000000";
				when "1111110011011" => data <= "000000";
				when "1111110011100" => data <= "000000";
				when "1111110011101" => data <= "000000";
				when "1111110011110" => data <= "000000";
				when "1111110011111" => data <= "000000";
				when "1111110100000" => data <= "000000";
				when "1111110100001" => data <= "000000";
				when "1111110100010" => data <= "000000";
				when "1111110100011" => data <= "000000";
				when "1111110100100" => data <= "000000";
				when "1111110100101" => data <= "000000";
				when "1111110100110" => data <= "000000";
				when "1111110100111" => data <= "000000";
				when "1111110101000" => data <= "000000";
				when "1111110101001" => data <= "000000";
				when "1111110101010" => data <= "100111";
				when "1111110101011" => data <= "100111";
				when "1111110101100" => data <= "010011";
				when "1111110101101" => data <= "010011";
				when "1111110101110" => data <= "100111";
				when "1111110101111" => data <= "100111";
				when "1111110110000" => data <= "000000";
				when "1111110110001" => data <= "000000";
				when "1111110110010" => data <= "000000";
				when "1111110110011" => data <= "000000";
				when "1111110110100" => data <= "000000";
				when "1111110110101" => data <= "000000";
				when "1111110110110" => data <= "000000";
				when "1111110110111" => data <= "010011";
				when "1111110111000" => data <= "111111";
				when "1111110111001" => data <= "010011";
				when "1111110111010" => data <= "010011";
				when "1111110111011" => data <= "010011";
				when "1111110111100" => data <= "010011";
				when "1111110111101" => data <= "000000";
				when "1111110111110" => data <= "000000";
				when "1111110111111" => data <= "000000";
				when "1111111000000" => data <= "010011";
				when "1111111000001" => data <= "111111";
				when "1111111000010" => data <= "010011";
				when "1111111000011" => data <= "010011";
				when "1111111000100" => data <= "010011";
				when "1111111000101" => data <= "010011";
				when "1111111000110" => data <= "000000";
				when "1111111000111" => data <= "000000";
				when "1111111001000" => data <= "000000";
				when "1111111001001" => data <= "000000";
				when "1111111001010" => data <= "000000";
				when "1111111001011" => data <= "100111";
				when "1111111001100" => data <= "100111";
				when "1111111001101" => data <= "010011";
				when "1111111001110" => data <= "010011";
				when "1111111001111" => data <= "010011";
				when "1111111010000" => data <= "100111";
				when "1111111010001" => data <= "100111";
				when "1111111010010" => data <= "000000";
				when "1111111010011" => data <= "000000";
				when "1111111010100" => data <= "000000";
				when "1111111010101" => data <= "000000";
				when "1111111010110" => data <= "000000";
				when "1111111010111" => data <= "000000";
				when "1111111011000" => data <= "000000";
				when "1111111011001" => data <= "000000";
				when "1111111011010" => data <= "000000";
				when "1111111011011" => data <= "000000";
				when "1111111011100" => data <= "000000";
				when "1111111011101" => data <= "000000";
				when "1111111011110" => data <= "000000";
				when "1111111011111" => data <= "000000";
				when "1111111100000" => data <= "000000";
				when "1111111100001" => data <= "000000";
				when "1111111100010" => data <= "000000";
				when "1111111100011" => data <= "000000";
				when "1111111100100" => data <= "000000";
				when "1111111100101" => data <= "000000";
				when "1111111100110" => data <= "000000";
				when "1111111100111" => data <= "000000";
				when "1111111101000" => data <= "000000";
				when "1111111101001" => data <= "000000";
				when "1111111101010" => data <= "000000";
				when "1111111101011" => data <= "000000";
				when "1111111101100" => data <= "000000";
				when "1111111101101" => data <= "000000";
				when "1111111101110" => data <= "000000";
				when "1111111101111" => data <= "000000";
				when "1111111110000" => data <= "000000";
				when "1111111110001" => data <= "000000";
				when "1111111110010" => data <= "000000";
				when "1111111110011" => data <= "000000";
				when "1111111110100" => data <= "000000";
				when "1111111110101" => data <= "000000";
				when "1111111110110" => data <= "000000";
				when "1111111110111" => data <= "000000";
				when "1111111111000" => data <= "000000";
				when "1111111111001" => data <= "000000";
				when "1111111111010" => data <= "000000";
				when "1111111111011" => data <= "000000";
				when "1111111111100" => data <= "000000";
				when "1111111111101" => data <= "000000";
				when "1111111111110" => data <= "000000";
				when "1111111111111" => data <= "000000";
				when "10000000000000" => data <= "000000";
				when "10000000000001" => data <= "000000";
				when "10000000000010" => data <= "000000";
				when "10000000000011" => data <= "000000";
				when "10000000000100" => data <= "000000";
				when "10000000000101" => data <= "000000";
				when "10000000000110" => data <= "000000";
				when "10000000000111" => data <= "000000";
				when "10000000001000" => data <= "000000";
				when "10000000001001" => data <= "000000";
				when "10000000001010" => data <= "000000";
				when "10000000001011" => data <= "000000";
				when "10000000001100" => data <= "000000";
				when "10000000001101" => data <= "000000";
				when "10000000001110" => data <= "000000";
				when "10000000001111" => data <= "000000";
				when "10000000010000" => data <= "000000";
				when "10000000010001" => data <= "000000";
				when "10000000010010" => data <= "000000";
				when "10000000010011" => data <= "000000";
				when "10000000010100" => data <= "000000";
				when "10000000010101" => data <= "000000";
				when "10000000010110" => data <= "000000";
				when "10000000010111" => data <= "000000";
				when "10000000011000" => data <= "000000";
				when "10000000011001" => data <= "000000";
				when "10000000011010" => data <= "000000";
				when "10000000011011" => data <= "000000";
				when "10000000011100" => data <= "000000";
				when "10000000011101" => data <= "000000";
				when "10000000011110" => data <= "000000";
				when "10000000011111" => data <= "000000";
				when "10000000100000" => data <= "000000";
				when "10000000100001" => data <= "000000";
				when "10000000100010" => data <= "000000";
				when "10000000100011" => data <= "000000";
				when "10000000100100" => data <= "000000";
				when "10000000100101" => data <= "000000";
				when "10000000100110" => data <= "000000";
				when "10000000100111" => data <= "000000";
				when "10000000101000" => data <= "000000";
				when "10000000101001" => data <= "000000";
				when "10000000101010" => data <= "100011";
				when "10000000101011" => data <= "100111";
				when "10000000101100" => data <= "100111";
				when "10000000101101" => data <= "100111";
				when "10000000101110" => data <= "100111";
				when "10000000101111" => data <= "100011";
				when "10000000110000" => data <= "000000";
				when "10000000110001" => data <= "000000";
				when "10000000110010" => data <= "000000";
				when "10000000110011" => data <= "000000";
				when "10000000110100" => data <= "000000";
				when "10000000110101" => data <= "000000";
				when "10000000110110" => data <= "000000";
				when "10000000110111" => data <= "100111";
				when "10000000111000" => data <= "100111";
				when "10000000111001" => data <= "010011";
				when "10000000111010" => data <= "010011";
				when "10000000111011" => data <= "100111";
				when "10000000111100" => data <= "100111";
				when "10000000111101" => data <= "000000";
				when "10000000111110" => data <= "000000";
				when "10000000111111" => data <= "000000";
				when "10000001000000" => data <= "100111";
				when "10000001000001" => data <= "100111";
				when "10000001000010" => data <= "010011";
				when "10000001000011" => data <= "010011";
				when "10000001000100" => data <= "100111";
				when "10000001000101" => data <= "100111";
				when "10000001000110" => data <= "000000";
				when "10000001000111" => data <= "000000";
				when "10000001001000" => data <= "000000";
				when "10000001001001" => data <= "000000";
				when "10000001001010" => data <= "000000";
				when "10000001001011" => data <= "100011";
				when "10000001001100" => data <= "100111";
				when "10000001001101" => data <= "100111";
				when "10000001001110" => data <= "010011";
				when "10000001001111" => data <= "100111";
				when "10000001010000" => data <= "100111";
				when "10000001010001" => data <= "100011";
				when "10000001010010" => data <= "000000";
				when "10000001010011" => data <= "000000";
				when "10000001010100" => data <= "000000";
				when "10000001010101" => data <= "000000";
				when "10000001010110" => data <= "000000";
				when "10000001010111" => data <= "000000";
				when "10000001011000" => data <= "000000";
				when "10000001011001" => data <= "000000";
				when "10000001011010" => data <= "000000";
				when "10000001011011" => data <= "000000";
				when "10000001011100" => data <= "000000";
				when "10000001011101" => data <= "000000";
				when "10000001011110" => data <= "000000";
				when "10000001011111" => data <= "000000";
				when "10000001100000" => data <= "000000";
				when "10000001100001" => data <= "000000";
				when "10000001100010" => data <= "000000";
				when "10000001100011" => data <= "000000";
				when "10000001100100" => data <= "000000";
				when "10000001100101" => data <= "000000";
				when "10000001100110" => data <= "000000";
				when "10000001100111" => data <= "000000";
				when "10000001101000" => data <= "000000";
				when "10000001101001" => data <= "000000";
				when "10000001101010" => data <= "000000";
				when "10000001101011" => data <= "000000";
				when "10000001101100" => data <= "000000";
				when "10000001101101" => data <= "000000";
				when "10000001101110" => data <= "000000";
				when "10000001101111" => data <= "000000";
				when "10000001110000" => data <= "000000";
				when "10000001110001" => data <= "000000";
				when "10000001110010" => data <= "000000";
				when "10000001110011" => data <= "000000";
				when "10000001110100" => data <= "000000";
				when "10000001110101" => data <= "000000";
				when "10000001110110" => data <= "000000";
				when "10000001110111" => data <= "000000";
				when "10000001111000" => data <= "000000";
				when "10000001111001" => data <= "000000";
				when "10000001111010" => data <= "000000";
				when "10000001111011" => data <= "000000";
				when "10000001111100" => data <= "000000";
				when "10000001111101" => data <= "000000";
				when "10000001111110" => data <= "000000";
				when "10000001111111" => data <= "000000";
				when "10000010000000" => data <= "000000";
				when "10000010000001" => data <= "000000";
				when "10000010000010" => data <= "000000";
				when "10000010000011" => data <= "000000";
				when "10000010000100" => data <= "000000";
				when "10000010000101" => data <= "000000";
				when "10000010000110" => data <= "000000";
				when "10000010000111" => data <= "000000";
				when "10000010001000" => data <= "000000";
				when "10000010001001" => data <= "000000";
				when "10000010001010" => data <= "000000";
				when "10000010001011" => data <= "000000";
				when "10000010001100" => data <= "000000";
				when "10000010001101" => data <= "000000";
				when "10000010001110" => data <= "000000";
				when "10000010001111" => data <= "000000";
				when "10000010010000" => data <= "000000";
				when "10000010010001" => data <= "000000";
				when "10000010010010" => data <= "000000";
				when "10000010010011" => data <= "000000";
				when "10000010010100" => data <= "000000";
				when "10000010010101" => data <= "000000";
				when "10000010010110" => data <= "000000";
				when "10000010010111" => data <= "000000";
				when "10000010011000" => data <= "000000";
				when "10000010011001" => data <= "000000";
				when "10000010011010" => data <= "000000";
				when "10000010011011" => data <= "000000";
				when "10000010011100" => data <= "000000";
				when "10000010011101" => data <= "000000";
				when "10000010011110" => data <= "000000";
				when "10000010011111" => data <= "000000";
				when "10000010100000" => data <= "000000";
				when "10000010100001" => data <= "000000";
				when "10000010100010" => data <= "000000";
				when "10000010100011" => data <= "000000";
				when "10000010100100" => data <= "000000";
				when "10000010100101" => data <= "000000";
				when "10000010100110" => data <= "000000";
				when "10000010100111" => data <= "000000";
				when "10000010101000" => data <= "000000";
				when "10000010101001" => data <= "000000";
				when "10000010101010" => data <= "100011";
				when "10000010101011" => data <= "100011";
				when "10000010101100" => data <= "100111";
				when "10000010101101" => data <= "100111";
				when "10000010101110" => data <= "100011";
				when "10000010101111" => data <= "100011";
				when "10000010110000" => data <= "000000";
				when "10000010110001" => data <= "000000";
				when "10000010110010" => data <= "000000";
				when "10000010110011" => data <= "000000";
				when "10000010110100" => data <= "000000";
				when "10000010110101" => data <= "000000";
				when "10000010110110" => data <= "000000";
				when "10000010110111" => data <= "100011";
				when "10000010111000" => data <= "100111";
				when "10000010111001" => data <= "100111";
				when "10000010111010" => data <= "100111";
				when "10000010111011" => data <= "100111";
				when "10000010111100" => data <= "100011";
				when "10000010111101" => data <= "000000";
				when "10000010111110" => data <= "000000";
				when "10000010111111" => data <= "000000";
				when "10000011000000" => data <= "100011";
				when "10000011000001" => data <= "100111";
				when "10000011000010" => data <= "100111";
				when "10000011000011" => data <= "100111";
				when "10000011000100" => data <= "100111";
				when "10000011000101" => data <= "100011";
				when "10000011000110" => data <= "000000";
				when "10000011000111" => data <= "000000";
				when "10000011001000" => data <= "000000";
				when "10000011001001" => data <= "000000";
				when "10000011001010" => data <= "000000";
				when "10000011001011" => data <= "100011";
				when "10000011001100" => data <= "100011";
				when "10000011001101" => data <= "100111";
				when "10000011001110" => data <= "100111";
				when "10000011001111" => data <= "100111";
				when "10000011010000" => data <= "100011";
				when "10000011010001" => data <= "100011";
				when "10000011010010" => data <= "000000";
				when "10000011010011" => data <= "000000";
				when "10000011010100" => data <= "000000";
				when "10000011010101" => data <= "000000";
				when "10000011010110" => data <= "000000";
				when "10000011010111" => data <= "000000";
				when "10000011011000" => data <= "000000";
				when "10000011011001" => data <= "000000";
				when "10000011011010" => data <= "000000";
				when "10000011011011" => data <= "000000";
				when "10000011011100" => data <= "000000";
				when "10000011011101" => data <= "000000";
				when "10000011011110" => data <= "000000";
				when "10000011011111" => data <= "000000";
				when "10000011100000" => data <= "000000";
				when "10000011100001" => data <= "000000";
				when "10000011100010" => data <= "000000";
				when "10000011100011" => data <= "000000";
				when "10000011100100" => data <= "000000";
				when "10000011100101" => data <= "000000";
				when "10000011100110" => data <= "000000";
				when "10000011100111" => data <= "000000";
				when "10000011101000" => data <= "000000";
				when "10000011101001" => data <= "000000";
				when "10000011101010" => data <= "000000";
				when "10000011101011" => data <= "000000";
				when "10000011101100" => data <= "000000";
				when "10000011101101" => data <= "000000";
				when "10000011101110" => data <= "000000";
				when "10000011101111" => data <= "000000";
				when "10000011110000" => data <= "000000";
				when "10000011110001" => data <= "000000";
				when "10000011110010" => data <= "000000";
				when "10000011110011" => data <= "000000";
				when "10000011110100" => data <= "000000";
				when "10000011110101" => data <= "000000";
				when "10000011110110" => data <= "000000";
				when "10000011110111" => data <= "000000";
				when "10000011111000" => data <= "000000";
				when "10000011111001" => data <= "000000";
				when "10000011111010" => data <= "000000";
				when "10000011111011" => data <= "000000";
				when "10000011111100" => data <= "000000";
				when "10000011111101" => data <= "000000";
				when "10000011111110" => data <= "000000";
				when "10000011111111" => data <= "000000";
				when "10000100000000" => data <= "000000";
				when "10000100000001" => data <= "000000";
				when "10000100000010" => data <= "000000";
				when "10000100000011" => data <= "000000";
				when "10000100000100" => data <= "000000";
				when "10000100000101" => data <= "000000";
				when "10000100000110" => data <= "000000";
				when "10000100000111" => data <= "000000";
				when "10000100001000" => data <= "000000";
				when "10000100001001" => data <= "000000";
				when "10000100001010" => data <= "000000";
				when "10000100001011" => data <= "000000";
				when "10000100001100" => data <= "000000";
				when "10000100001101" => data <= "000000";
				when "10000100001110" => data <= "000000";
				when "10000100001111" => data <= "000000";
				when "10000100010000" => data <= "000000";
				when "10000100010001" => data <= "000000";
				when "10000100010010" => data <= "000000";
				when "10000100010011" => data <= "000000";
				when "10000100010100" => data <= "000000";
				when "10000100010101" => data <= "000000";
				when "10000100010110" => data <= "000000";
				when "10000100010111" => data <= "000000";
				when "10000100011000" => data <= "000000";
				when "10000100011001" => data <= "000000";
				when "10000100011010" => data <= "000000";
				when "10000100011011" => data <= "000000";
				when "10000100011100" => data <= "000000";
				when "10000100011101" => data <= "000000";
				when "10000100011110" => data <= "000000";
				when "10000100011111" => data <= "000000";
				when "10000100100000" => data <= "000000";
				when "10000100100001" => data <= "000000";
				when "10000100100010" => data <= "000000";
				when "10000100100011" => data <= "000000";
				when "10000100100100" => data <= "000000";
				when "10000100100101" => data <= "000000";
				when "10000100100110" => data <= "000000";
				when "10000100100111" => data <= "000000";
				when "10000100101000" => data <= "000000";
				when "10000100101001" => data <= "000000";
				when "10000100101010" => data <= "000000";
				when "10000100101011" => data <= "100011";
				when "10000100101100" => data <= "100011";
				when "10000100101101" => data <= "100011";
				when "10000100101110" => data <= "100011";
				when "10000100101111" => data <= "000000";
				when "10000100110000" => data <= "000000";
				when "10000100110001" => data <= "000000";
				when "10000100110010" => data <= "000000";
				when "10000100110011" => data <= "000000";
				when "10000100110100" => data <= "000000";
				when "10000100110101" => data <= "000000";
				when "10000100110110" => data <= "000000";
				when "10000100110111" => data <= "100011";
				when "10000100111000" => data <= "100011";
				when "10000100111001" => data <= "100111";
				when "10000100111010" => data <= "100111";
				when "10000100111011" => data <= "100011";
				when "10000100111100" => data <= "100011";
				when "10000100111101" => data <= "000000";
				when "10000100111110" => data <= "000000";
				when "10000100111111" => data <= "000000";
				when "10000101000000" => data <= "100011";
				when "10000101000001" => data <= "100011";
				when "10000101000010" => data <= "100111";
				when "10000101000011" => data <= "100111";
				when "10000101000100" => data <= "100011";
				when "10000101000101" => data <= "100011";
				when "10000101000110" => data <= "000000";
				when "10000101000111" => data <= "000000";
				when "10000101001000" => data <= "000000";
				when "10000101001001" => data <= "000000";
				when "10000101001010" => data <= "000000";
				when "10000101001011" => data <= "000000";
				when "10000101001100" => data <= "100011";
				when "10000101001101" => data <= "100011";
				when "10000101001110" => data <= "100011";
				when "10000101001111" => data <= "100011";
				when "10000101010000" => data <= "100011";
				when "10000101010001" => data <= "000000";
				when "10000101010010" => data <= "000000";
				when "10000101010011" => data <= "000000";
				when "10000101010100" => data <= "000000";
				when "10000101010101" => data <= "000000";
				when "10000101010110" => data <= "000000";
				when "10000101010111" => data <= "000000";
				when "10000101011000" => data <= "000000";
				when "10000101011001" => data <= "000000";
				when "10000101011010" => data <= "000000";
				when "10000101011011" => data <= "000000";
				when "10000101011100" => data <= "000000";
				when "10000101011101" => data <= "000000";
				when "10000101011110" => data <= "000000";
				when "10000101011111" => data <= "000000";
				when "10000101100000" => data <= "000000";
				when "10000101100001" => data <= "000000";
				when "10000101100010" => data <= "000000";
				when "10000101100011" => data <= "000000";
				when "10000101100100" => data <= "000000";
				when "10000101100101" => data <= "000000";
				when "10000101100110" => data <= "000000";
				when "10000101100111" => data <= "000000";
				when "10000101101000" => data <= "000000";
				when "10000101101001" => data <= "000000";
				when "10000101101010" => data <= "000000";
				when "10000101101011" => data <= "000000";
				when "10000101101100" => data <= "000000";
				when "10000101101101" => data <= "000000";
				when "10000101101110" => data <= "000000";
				when "10000101101111" => data <= "000000";
				when "10000101110000" => data <= "000000";
				when "10000101110001" => data <= "000000";
				when "10000101110010" => data <= "000000";
				when "10000101110011" => data <= "000000";
				when "10000101110100" => data <= "000000";
				when "10000101110101" => data <= "000000";
				when "10000101110110" => data <= "000000";
				when "10000101110111" => data <= "000000";
				when "10000101111000" => data <= "000000";
				when "10000101111001" => data <= "000000";
				when "10000101111010" => data <= "000000";
				when "10000101111011" => data <= "000000";
				when "10000101111100" => data <= "000000";
				when "10000101111101" => data <= "000000";
				when "10000101111110" => data <= "000000";
				when "10000101111111" => data <= "000000";
				when "10000110000000" => data <= "000000";
				when "10000110000001" => data <= "000000";
				when "10000110000010" => data <= "000000";
				when "10000110000011" => data <= "000000";
				when "10000110000100" => data <= "000000";
				when "10000110000101" => data <= "000000";
				when "10000110000110" => data <= "000000";
				when "10000110000111" => data <= "000000";
				when "10000110001000" => data <= "000000";
				when "10000110001001" => data <= "000000";
				when "10000110001010" => data <= "000000";
				when "10000110001011" => data <= "000000";
				when "10000110001100" => data <= "000000";
				when "10000110001101" => data <= "000000";
				when "10000110001110" => data <= "000000";
				when "10000110001111" => data <= "000000";
				when "10000110010000" => data <= "000000";
				when "10000110010001" => data <= "000000";
				when "10000110010010" => data <= "000000";
				when "10000110010011" => data <= "000000";
				when "10000110010100" => data <= "000000";
				when "10000110010101" => data <= "000000";
				when "10000110010110" => data <= "000000";
				when "10000110010111" => data <= "000000";
				when "10000110011000" => data <= "000000";
				when "10000110011001" => data <= "000000";
				when "10000110011010" => data <= "000000";
				when "10000110011011" => data <= "000000";
				when "10000110011100" => data <= "000000";
				when "10000110011101" => data <= "000000";
				when "10000110011110" => data <= "000000";
				when "10000110011111" => data <= "000000";
				when "10000110100000" => data <= "000000";
				when "10000110100001" => data <= "000000";
				when "10000110100010" => data <= "000000";
				when "10000110100011" => data <= "000000";
				when "10000110100100" => data <= "000000";
				when "10000110100101" => data <= "000000";
				when "10000110100110" => data <= "000000";
				when "10000110100111" => data <= "000000";
				when "10000110101000" => data <= "000000";
				when "10000110101001" => data <= "000000";
				when "10000110101010" => data <= "000000";
				when "10000110101011" => data <= "000000";
				when "10000110101100" => data <= "000000";
				when "10000110101101" => data <= "000000";
				when "10000110101110" => data <= "000000";
				when "10000110101111" => data <= "000000";
				when "10000110110000" => data <= "000000";
				when "10000110110001" => data <= "000000";
				when "10000110110010" => data <= "000000";
				when "10000110110011" => data <= "000000";
				when "10000110110100" => data <= "000000";
				when "10000110110101" => data <= "000000";
				when "10000110110110" => data <= "000000";
				when "10000110110111" => data <= "000000";
				when "10000110111000" => data <= "100011";
				when "10000110111001" => data <= "100011";
				when "10000110111010" => data <= "100011";
				when "10000110111011" => data <= "100011";
				when "10000110111100" => data <= "000000";
				when "10000110111101" => data <= "000000";
				when "10000110111110" => data <= "000000";
				when "10000110111111" => data <= "000000";
				when "10000111000000" => data <= "000000";
				when "10000111000001" => data <= "100011";
				when "10000111000010" => data <= "100011";
				when "10000111000011" => data <= "100011";
				when "10000111000100" => data <= "100011";
				when "10000111000101" => data <= "000000";
				when "10000111000110" => data <= "000000";
				when "10000111000111" => data <= "000000";
				when "10000111001000" => data <= "000000";
				when "10000111001001" => data <= "000000";
				when "10000111001010" => data <= "000000";
				when "10000111001011" => data <= "000000";
				when "10000111001100" => data <= "000000";
				when "10000111001101" => data <= "000000";
				when "10000111001110" => data <= "000000";
				when "10000111001111" => data <= "000000";
				when "10000111010000" => data <= "000000";
				when "10000111010001" => data <= "000000";
				when "10000111010010" => data <= "000000";
				when "10000111010011" => data <= "000000";
				when "10000111010100" => data <= "000000";
				when "10000111010101" => data <= "000000";
				when "10000111010110" => data <= "000000";
				when "10000111010111" => data <= "000000";
				when "10000111011000" => data <= "000000";
				when "10000111011001" => data <= "000000";
				when "10000111011010" => data <= "000000";
				when "10000111011011" => data <= "000000";
				when "10000111011100" => data <= "000000";
				when "10000111011101" => data <= "000000";
				when "10000111011110" => data <= "000000";
				when "10000111011111" => data <= "000000";
				when "10000111100000" => data <= "000000";
				when "10000111100001" => data <= "000000";
				when "10000111100010" => data <= "000000";
				when "10000111100011" => data <= "000000";
				when "10000111100100" => data <= "000000";
				when "10000111100101" => data <= "000000";
				when "10000111100110" => data <= "000000";
				when "10000111100111" => data <= "000000";
				when "10000111101000" => data <= "000000";
				when "10000111101001" => data <= "000000";
				when "10000111101010" => data <= "000000";
				when "10000111101011" => data <= "000000";
				when "10000111101100" => data <= "000000";
				when "10000111101101" => data <= "000000";
				when "10000111101110" => data <= "000000";
				when "10000111101111" => data <= "000000";
				when "10000111110000" => data <= "000000";
				when "10000111110001" => data <= "000000";
				when "10000111110010" => data <= "000000";
				when "10000111110011" => data <= "000000";
				when "10000111110100" => data <= "000000";
				when "10000111110101" => data <= "000000";
				when "10000111110110" => data <= "000000";
				when "10000111110111" => data <= "000000";
				when "10000111111000" => data <= "000000";
				when "10000111111001" => data <= "000000";
				when "10000111111010" => data <= "000000";
				when "10000111111011" => data <= "000000";
				when "10000111111100" => data <= "000000";
				when "10000111111101" => data <= "000000";
				when "10000111111110" => data <= "000000";
				when "10000111111111" => data <= "000000";
				when "10001000000000" => data <= "000000";
				when "10001000000001" => data <= "000000";
				when "10001000000010" => data <= "000000";
				when "10001000000011" => data <= "000000";
				when "10001000000100" => data <= "000000";
				when "10001000000101" => data <= "000000";
				when "10001000000110" => data <= "000000";
				when "10001000000111" => data <= "000000";
				when "10001000001000" => data <= "000000";
				when "10001000001001" => data <= "000000";
				when "10001000001010" => data <= "000000";
				when "10001000001011" => data <= "000000";
				when "10001000001100" => data <= "000000";
				when "10001000001101" => data <= "000000";
				when "10001000001110" => data <= "000000";
				when "10001000001111" => data <= "000000";
				when "10001000010000" => data <= "000000";
				when "10001000010001" => data <= "000000";
				when "10001000010010" => data <= "000000";
				when "10001000010011" => data <= "000000";
				when "10001000010100" => data <= "000000";
				when "10001000010101" => data <= "000000";
				when "10001000010110" => data <= "000000";
				when "10001000010111" => data <= "000000";
				when "10001000011000" => data <= "000000";
				when "10001000011001" => data <= "000000";
				when "10001000011010" => data <= "000000";
				when "10001000011011" => data <= "000000";
				when "10001000011100" => data <= "000000";
				when "10001000011101" => data <= "000000";
				when "10001000011110" => data <= "000000";
				when "10001000011111" => data <= "000000";
				when "10001000100000" => data <= "000000";
				when "10001000100001" => data <= "000000";
				when "10001000100010" => data <= "000000";
				when "10001000100011" => data <= "000000";
				when "10001000100100" => data <= "000000";
				when "10001000100101" => data <= "000000";
				when "10001000100110" => data <= "000000";
				when "10001000100111" => data <= "000000";
				when "10001000101000" => data <= "000000";
				when "10001000101001" => data <= "000000";
				when "10001000101010" => data <= "000000";
				when "10001000101011" => data <= "000000";
				when "10001000101100" => data <= "000000";
				when "10001000101101" => data <= "000000";
				when "10001000101110" => data <= "000000";
				when "10001000101111" => data <= "000000";
				when "10001000110000" => data <= "000000";
				when "10001000110001" => data <= "000000";
				when "10001000110010" => data <= "000000";
				when "10001000110011" => data <= "000000";
				when "10001000110100" => data <= "000000";
				when "10001000110101" => data <= "000000";
				when "10001000110110" => data <= "000000";
				when "10001000110111" => data <= "000000";
				when "10001000111000" => data <= "000000";
				when "10001000111001" => data <= "000000";
				when "10001000111010" => data <= "000000";
				when "10001000111011" => data <= "000000";
				when "10001000111100" => data <= "000000";
				when "10001000111101" => data <= "000000";
				when "10001000111110" => data <= "000000";
				when "10001000111111" => data <= "000000";
				when "10001001000000" => data <= "000000";
				when "10001001000001" => data <= "000000";
				when "10001001000010" => data <= "000000";
				when "10001001000011" => data <= "000000";
				when "10001001000100" => data <= "000000";
				when "10001001000101" => data <= "000000";
				when "10001001000110" => data <= "000000";
				when "10001001000111" => data <= "000000";
				when "10001001001000" => data <= "000000";
				when "10001001001001" => data <= "000000";
				when "10001001001010" => data <= "000000";
				when "10001001001011" => data <= "000000";
				when "10001001001100" => data <= "000000";
				when "10001001001101" => data <= "000000";
				when "10001001001110" => data <= "000000";
				when "10001001001111" => data <= "000000";
				when "10001001010000" => data <= "000000";
				when "10001001010001" => data <= "000000";
				when "10001001010010" => data <= "000000";
				when "10001001010011" => data <= "000000";
				when "10001001010100" => data <= "000000";
				when "10001001010101" => data <= "000000";
				when "10001001010110" => data <= "000000";
				when "10001001010111" => data <= "000000";
				when "10001001011000" => data <= "000000";
				when "10001001011001" => data <= "000000";
				when "10001001011010" => data <= "000000";
				when "10001001011011" => data <= "000000";
				when "10001001011100" => data <= "000000";
				when "10001001011101" => data <= "000000";
				when "10001001011110" => data <= "000000";
				when "10001001011111" => data <= "000000";
				when "10001001100000" => data <= "000000";
				when "10001001100001" => data <= "000000";
				when "10001001100010" => data <= "000000";
				when "10001001100011" => data <= "000000";
				when "10001001100100" => data <= "000000";
				when "10001001100101" => data <= "000000";
				when "10001001100110" => data <= "000000";
				when "10001001100111" => data <= "000000";
				when "10001001101000" => data <= "000000";
				when "10001001101001" => data <= "000000";
				when "10001001101010" => data <= "000000";
				when "10001001101011" => data <= "000000";
				when "10001001101100" => data <= "000000";
				when "10001001101101" => data <= "000000";
				when "10001001101110" => data <= "000000";
				when "10001001101111" => data <= "000000";
				when "10001001110000" => data <= "000000";
				when "10001001110001" => data <= "000000";
				when "10001001110010" => data <= "000000";
				when "10001001110011" => data <= "000000";
				when "10001001110100" => data <= "000000";
				when "10001001110101" => data <= "000000";
				when "10001001110110" => data <= "000000";
				when "10001001110111" => data <= "000000";
				when "10001001111000" => data <= "000000";
				when "10001001111001" => data <= "000000";
				when "10001001111010" => data <= "000000";
				when "10001001111011" => data <= "000000";
				when "10001001111100" => data <= "000000";
				when "10001001111101" => data <= "000000";
				when "10001001111110" => data <= "000000";
				when "10001001111111" => data <= "000000";
				when "10001010000000" => data <= "000000";
				when "10001010000001" => data <= "000000";
				when "10001010000010" => data <= "000000";
				when "10001010000011" => data <= "000000";
				when "10001010000100" => data <= "000000";
				when "10001010000101" => data <= "000000";
				when "10001010000110" => data <= "000000";
				when "10001010000111" => data <= "000000";
				when "10001010001000" => data <= "000000";
				when "10001010001001" => data <= "000000";
				when "10001010001010" => data <= "000000";
				when "10001010001011" => data <= "000000";
				when "10001010001100" => data <= "000000";
				when "10001010001101" => data <= "000000";
				when "10001010001110" => data <= "000000";
				when "10001010001111" => data <= "000000";
				when "10001010010000" => data <= "000000";
				when "10001010010001" => data <= "000000";
				when "10001010010010" => data <= "000000";
				when "10001010010011" => data <= "000000";
				when "10001010010100" => data <= "000000";
				when "10001010010101" => data <= "000000";
				when "10001010010110" => data <= "000000";
				when "10001010010111" => data <= "000000";
				when "10001010011000" => data <= "000000";
				when "10001010011001" => data <= "000000";
				when "10001010011010" => data <= "000000";
				when "10001010011011" => data <= "000000";
				when "10001010011100" => data <= "000000";
				when "10001010011101" => data <= "000000";
				when "10001010011110" => data <= "000000";
				when "10001010011111" => data <= "000000";
				when "10001010100000" => data <= "000000";
				when "10001010100001" => data <= "000000";
				when "10001010100010" => data <= "000000";
				when "10001010100011" => data <= "000000";
				when "10001010100100" => data <= "000000";
				when "10001010100101" => data <= "000000";
				when "10001010100110" => data <= "000000";
				when "10001010100111" => data <= "000000";
				when "10001010101000" => data <= "000000";
				when "10001010101001" => data <= "000000";
				when "10001010101010" => data <= "000000";
				when "10001010101011" => data <= "000000";
				when "10001010101100" => data <= "000000";
				when "10001010101101" => data <= "000000";
				when "10001010101110" => data <= "000000";
				when "10001010101111" => data <= "000000";
				when "10001010110000" => data <= "000000";
				when "10001010110001" => data <= "000000";
				when "10001010110010" => data <= "000000";
				when "10001010110011" => data <= "000000";
				when "10001010110100" => data <= "000000";
				when "10001010110101" => data <= "000000";
				when "10001010110110" => data <= "000000";
				when "10001010110111" => data <= "000000";
				when "10001010111000" => data <= "000000";
				when "10001010111001" => data <= "000000";
				when "10001010111010" => data <= "000000";
				when "10001010111011" => data <= "000000";
				when "10001010111100" => data <= "000000";
				when "10001010111101" => data <= "000000";
				when "10001010111110" => data <= "000000";
				when "10001010111111" => data <= "000000";
				when "10001011000000" => data <= "000000";
				when "10001011000001" => data <= "000000";
				when "10001011000010" => data <= "000000";
				when "10001011000011" => data <= "000000";
				when "10001011000100" => data <= "000000";
				when "10001011000101" => data <= "000000";
				when "10001011000110" => data <= "000000";
				when "10001011000111" => data <= "000000";
				when "10001011001000" => data <= "000000";
				when "10001011001001" => data <= "000000";
				when "10001011001010" => data <= "000000";
				when "10001011001011" => data <= "000000";
				when "10001011001100" => data <= "000000";
				when "10001011001101" => data <= "000000";
				when "10001011001110" => data <= "000000";
				when "10001011001111" => data <= "000000";
				when "10001011010000" => data <= "000000";
				when "10001011010001" => data <= "000000";
				when "10001011010010" => data <= "000000";
				when "10001011010011" => data <= "000000";
				when "10001011010100" => data <= "000000";
				when "10001011010101" => data <= "000000";
				when "10001011010110" => data <= "000000";
				when "10001011010111" => data <= "000000";
				when "10001011011000" => data <= "000000";
				when "10001011011001" => data <= "000000";
				when "10001011011010" => data <= "000000";
				when "10001011011011" => data <= "000000";
				when "10001011011100" => data <= "000000";
				when "10001011011101" => data <= "000000";
				when "10001011011110" => data <= "000000";
				when "10001011011111" => data <= "000000";
				when "10001011100000" => data <= "000000";
				when "10001011100001" => data <= "000000";
				when "10001011100010" => data <= "000000";
				when "10001011100011" => data <= "000000";
				when "10001011100100" => data <= "000000";
				when "10001011100101" => data <= "000000";
				when "10001011100110" => data <= "000000";
				when "10001011100111" => data <= "000000";
				when "10001011101000" => data <= "000000";
				when "10001011101001" => data <= "000000";
				when "10001011101010" => data <= "000000";
				when "10001011101011" => data <= "000000";
				when "10001011101100" => data <= "000000";
				when "10001011101101" => data <= "000000";
				when "10001011101110" => data <= "000000";
				when "10001011101111" => data <= "000000";
				when "10001011110000" => data <= "000000";
				when "10001011110001" => data <= "000000";
				when "10001011110010" => data <= "000000";
				when "10001011110011" => data <= "000000";
				when "10001011110100" => data <= "000000";
				when "10001011110101" => data <= "000000";
				when "10001011110110" => data <= "000000";
				when "10001011110111" => data <= "000000";
				when "10001011111000" => data <= "000000";
				when "10001011111001" => data <= "000000";
				when "10001011111010" => data <= "000000";
				when "10001011111011" => data <= "000000";
				when "10001011111100" => data <= "000000";
				when "10001011111101" => data <= "000000";
				when "10001011111110" => data <= "000000";
				when "10001011111111" => data <= "000000";
				when "10001100000000" => data <= "000000";
				when "10001100000001" => data <= "000000";
				when "10001100000010" => data <= "000000";
				when "10001100000011" => data <= "000000";
				when "10001100000100" => data <= "000000";
				when "10001100000101" => data <= "000000";
				when "10001100000110" => data <= "000000";
				when "10001100000111" => data <= "000000";
				when "10001100001000" => data <= "000000";
				when "10001100001001" => data <= "000000";
				when "10001100001010" => data <= "000000";
				when "10001100001011" => data <= "000000";
				when "10001100001100" => data <= "000000";
				when "10001100001101" => data <= "000000";
				when "10001100001110" => data <= "000000";
				when "10001100001111" => data <= "000000";
				when "10001100010000" => data <= "000000";
				when "10001100010001" => data <= "000000";
				when "10001100010010" => data <= "000000";
				when "10001100010011" => data <= "000000";
				when "10001100010100" => data <= "000000";
				when "10001100010101" => data <= "000000";
				when "10001100010110" => data <= "000000";
				when "10001100010111" => data <= "000000";
				when "10001100011000" => data <= "000000";
				when "10001100011001" => data <= "000000";
				when "10001100011010" => data <= "000000";
				when "10001100011011" => data <= "000000";
				when "10001100011100" => data <= "000000";
				when "10001100011101" => data <= "000000";
				when "10001100011110" => data <= "000000";
				when "10001100011111" => data <= "000000";
				when "10001100100000" => data <= "000000";
				when "10001100100001" => data <= "000000";
				when "10001100100010" => data <= "000000";
				when "10001100100011" => data <= "000000";
				when "10001100100100" => data <= "000000";
				when "10001100100101" => data <= "000000";
				when "10001100100110" => data <= "000000";
				when "10001100100111" => data <= "000000";
				when "10001100101000" => data <= "000000";
				when "10001100101001" => data <= "000000";
				when "10001100101010" => data <= "000000";
				when "10001100101011" => data <= "000000";
				when "10001100101100" => data <= "000000";
				when "10001100101101" => data <= "000000";
				when "10001100101110" => data <= "000000";
				when "10001100101111" => data <= "000000";
				when "10001100110000" => data <= "000000";
				when "10001100110001" => data <= "000000";
				when "10001100110010" => data <= "000000";
				when "10001100110011" => data <= "000000";
				when "10001100110100" => data <= "000000";
				when "10001100110101" => data <= "000000";
				when "10001100110110" => data <= "000000";
				when "10001100110111" => data <= "000000";
				when "10001100111000" => data <= "000000";
				when "10001100111001" => data <= "000000";
				when "10001100111010" => data <= "000000";
				when "10001100111011" => data <= "000000";
				when "10001100111100" => data <= "000000";
				when "10001100111101" => data <= "000000";
				when "10001100111110" => data <= "000000";
				when "10001100111111" => data <= "000000";
				when "10001101000000" => data <= "000000";
				when "10001101000001" => data <= "000000";
				when "10001101000010" => data <= "000000";
				when "10001101000011" => data <= "000000";
				when "10001101000100" => data <= "000000";
				when "10001101000101" => data <= "000000";
				when "10001101000110" => data <= "000000";
				when "10001101000111" => data <= "000000";
				when "10001101001000" => data <= "000000";
				when "10001101001001" => data <= "000000";
				when "10001101001010" => data <= "000000";
				when "10001101001011" => data <= "000000";
				when "10001101001100" => data <= "000000";
				when "10001101001101" => data <= "000000";
				when "10001101001110" => data <= "000000";
				when "10001101001111" => data <= "000000";
				when "10001101010000" => data <= "000000";
				when "10001101010001" => data <= "000000";
				when "10001101010010" => data <= "000000";
				when "10001101010011" => data <= "000000";
				when "10001101010100" => data <= "000000";
				when "10001101010101" => data <= "000000";
				when "10001101010110" => data <= "000000";
				when "10001101010111" => data <= "000000";
				when "10001101011000" => data <= "000000";
				when "10001101011001" => data <= "000000";
				when "10001101011010" => data <= "000000";
				when "10001101011011" => data <= "000000";
				when "10001101011100" => data <= "000000";
				when "10001101011101" => data <= "000000";
				when "10001101011110" => data <= "000000";
				when "10001101011111" => data <= "000000";
				when "10001101100000" => data <= "000000";
				when "10001101100001" => data <= "000000";
				when "10001101100010" => data <= "000000";
				when "10001101100011" => data <= "000000";
				when "10001101100100" => data <= "000000";
				when "10001101100101" => data <= "000000";
				when "10001101100110" => data <= "000000";
				when "10001101100111" => data <= "000000";
				when "10001101101000" => data <= "000000";
				when "10001101101001" => data <= "000000";
				when "10001101101010" => data <= "000000";
				when "10001101101011" => data <= "000000";
				when "10001101101100" => data <= "000000";
				when "10001101101101" => data <= "000000";
				when "10001101101110" => data <= "000000";
				when "10001101101111" => data <= "000000";
				when "10001101110000" => data <= "000000";
				when "10001101110001" => data <= "000000";
				when "10001101110010" => data <= "000000";
				when "10001101110011" => data <= "000000";
				when "10001101110100" => data <= "000000";
				when "10001101110101" => data <= "000000";
				when "10001101110110" => data <= "000000";
				when "10001101110111" => data <= "000000";
				when "10001101111000" => data <= "000000";
				when "10001101111001" => data <= "000000";
				when "10001101111010" => data <= "000000";
				when "10001101111011" => data <= "000000";
				when "10001101111100" => data <= "000000";
				when "10001101111101" => data <= "000000";
				when "10001101111110" => data <= "000000";
				when "10001101111111" => data <= "000000";
				when "10001110000000" => data <= "000000";
				when "10001110000001" => data <= "000000";
				when "10001110000010" => data <= "000000";
				when "10001110000011" => data <= "000000";
				when "10001110000100" => data <= "000000";
				when "10001110000101" => data <= "000000";
				when "10001110000110" => data <= "000000";
				when "10001110000111" => data <= "000000";
				when "10001110001000" => data <= "000000";
				when "10001110001001" => data <= "000000";
				when "10001110001010" => data <= "000000";
				when "10001110001011" => data <= "000000";
				when "10001110001100" => data <= "000000";
				when "10001110001101" => data <= "000000";
				when "10001110001110" => data <= "000000";
				when "10001110001111" => data <= "000000";
				when "10001110010000" => data <= "000000";
				when "10001110010001" => data <= "000000";
				when "10001110010010" => data <= "000000";
				when "10001110010011" => data <= "000000";
				when "10001110010100" => data <= "000000";
				when "10001110010101" => data <= "000000";
				when "10001110010110" => data <= "000000";
				when "10001110010111" => data <= "000000";
				when "10001110011000" => data <= "000000";
				when "10001110011001" => data <= "000000";
				when "10001110011010" => data <= "000000";
				when "10001110011011" => data <= "000000";
				when "10001110011100" => data <= "000000";
				when "10001110011101" => data <= "000000";
				when "10001110011110" => data <= "000000";
				when "10001110011111" => data <= "000000";
				when "10001110100000" => data <= "000000";
				when "10001110100001" => data <= "000000";
				when "10001110100010" => data <= "000000";
				when "10001110100011" => data <= "000000";
				when "10001110100100" => data <= "000000";
				when "10001110100101" => data <= "000000";
				when "10001110100110" => data <= "000000";
				when "10001110100111" => data <= "000000";
				when "10001110101000" => data <= "000000";
				when "10001110101001" => data <= "000000";
				when "10001110101010" => data <= "000000";
				when "10001110101011" => data <= "000000";
				when "10001110101100" => data <= "000000";
				when "10001110101101" => data <= "000000";
				when "10001110101110" => data <= "000000";
				when "10001110101111" => data <= "000000";
				when "10001110110000" => data <= "000000";
				when "10001110110001" => data <= "000000";
				when "10001110110010" => data <= "000000";
				when "10001110110011" => data <= "000000";
				when "10001110110100" => data <= "000000";
				when "10001110110101" => data <= "000000";
				when "10001110110110" => data <= "000000";
				when "10001110110111" => data <= "000000";
				when "10001110111000" => data <= "000000";
				when "10001110111001" => data <= "000000";
				when "10001110111010" => data <= "000000";
				when "10001110111011" => data <= "000000";
				when "10001110111100" => data <= "000000";
				when "10001110111101" => data <= "000000";
				when "10001110111110" => data <= "000000";
				when "10001110111111" => data <= "000000";
				when "10001111000000" => data <= "000000";
				when "10001111000001" => data <= "000000";
				when "10001111000010" => data <= "000000";
				when "10001111000011" => data <= "000000";
				when "10001111000100" => data <= "000000";
				when "10001111000101" => data <= "000000";
				when "10001111000110" => data <= "000000";
				when "10001111000111" => data <= "000000";
				when "10001111001000" => data <= "000000";
				when "10001111001001" => data <= "000000";
				when "10001111001010" => data <= "000000";
				when "10001111001011" => data <= "000000";
				when "10001111001100" => data <= "000000";
				when "10001111001101" => data <= "000000";
				when "10001111001110" => data <= "000000";
				when "10001111001111" => data <= "000000";
				when "10001111010000" => data <= "000000";
				when "10001111010001" => data <= "000000";
				when "10001111010010" => data <= "000000";
				when "10001111010011" => data <= "000000";
				when "10001111010100" => data <= "000000";
				when "10001111010101" => data <= "000000";
				when "10001111010110" => data <= "000000";
				when "10001111010111" => data <= "000000";
				when "10001111011000" => data <= "000000";
				when "10001111011001" => data <= "000000";
				when "10001111011010" => data <= "000000";
				when "10001111011011" => data <= "000000";
				when "10001111011100" => data <= "000000";
				when "10001111011101" => data <= "000000";
				when "10001111011110" => data <= "000000";
				when "10001111011111" => data <= "000000";
				when "10001111100000" => data <= "000000";
				when "10001111100001" => data <= "000000";
				when "10001111100010" => data <= "000000";
				when "10001111100011" => data <= "000000";
				when "10001111100100" => data <= "000000";
				when "10001111100101" => data <= "000000";
				when "10001111100110" => data <= "000000";
				when "10001111100111" => data <= "000000";
				when "10001111101000" => data <= "000000";
				when "10001111101001" => data <= "000000";
				when "10001111101010" => data <= "000000";
				when "10001111101011" => data <= "000000";
				when "10001111101100" => data <= "000000";
				when "10001111101101" => data <= "000000";
				when "10001111101110" => data <= "000000";
				when "10001111101111" => data <= "000000";
				when "10001111110000" => data <= "000000";
				when "10001111110001" => data <= "000000";
				when "10001111110010" => data <= "000000";
				when "10001111110011" => data <= "000000";
				when "10001111110100" => data <= "000000";
				when "10001111110101" => data <= "000000";
				when "10001111110110" => data <= "000000";
				when "10001111110111" => data <= "000000";
				when "10001111111000" => data <= "000000";
				when "10001111111001" => data <= "000000";
				when "10001111111010" => data <= "000000";
				when "10001111111011" => data <= "000000";
				when "10001111111100" => data <= "000000";
				when "10001111111101" => data <= "000000";
				when "10001111111110" => data <= "000000";
				when "10001111111111" => data <= "000000";
				when "10010000000000" => data <= "000000";
				when "10010000000001" => data <= "000000";
				when "10010000000010" => data <= "000000";
				when "10010000000011" => data <= "000000";
				when "10010000000100" => data <= "000000";
				when "10010000000101" => data <= "000000";
				when "10010000000110" => data <= "000000";
				when "10010000000111" => data <= "000000";
				when "10010000001000" => data <= "000000";
				when "10010000001001" => data <= "000000";
				when "10010000001010" => data <= "000000";
				when "10010000001011" => data <= "000000";
				when "10010000001100" => data <= "000000";
				when "10010000001101" => data <= "000000";
				when "10010000001110" => data <= "000000";
				when "10010000001111" => data <= "000000";
				when "10010000010000" => data <= "000000";
				when "10010000010001" => data <= "000000";
				when "10010000010010" => data <= "000000";
				when "10010000010011" => data <= "000000";
				when "10010000010100" => data <= "000000";
				when "10010000010101" => data <= "000000";
				when "10010000010110" => data <= "000000";
				when "10010000010111" => data <= "000000";
				when "10010000011000" => data <= "000000";
				when "10010000011001" => data <= "000000";
				when "10010000011010" => data <= "000000";
				when "10010000011011" => data <= "000000";
				when "10010000011100" => data <= "000000";
				when "10010000011101" => data <= "000000";
				when "10010000011110" => data <= "000000";
				when "10010000011111" => data <= "000000";
				when "10010000100000" => data <= "000000";
				when "10010000100001" => data <= "000000";
				when "10010000100010" => data <= "000000";
				when "10010000100011" => data <= "000000";
				when "10010000100100" => data <= "000000";
				when "10010000100101" => data <= "000000";
				when "10010000100110" => data <= "000000";
				when "10010000100111" => data <= "000000";
				when "10010000101000" => data <= "000000";
				when "10010000101001" => data <= "000000";
				when "10010000101010" => data <= "000000";
				when "10010000101011" => data <= "000000";
				when "10010000101100" => data <= "000000";
				when "10010000101101" => data <= "000000";
				when "10010000101110" => data <= "000000";
				when "10010000101111" => data <= "000000";
				when "10010000110000" => data <= "000000";
				when "10010000110001" => data <= "000000";
				when "10010000110010" => data <= "000000";
				when "10010000110011" => data <= "000000";
				when "10010000110100" => data <= "000000";
				when "10010000110101" => data <= "000000";
				when "10010000110110" => data <= "000000";
				when "10010000110111" => data <= "000000";
				when "10010000111000" => data <= "000000";
				when "10010000111001" => data <= "000000";
				when "10010000111010" => data <= "000000";
				when "10010000111011" => data <= "000000";
				when "10010000111100" => data <= "000000";
				when "10010000111101" => data <= "000000";
				when "10010000111110" => data <= "000000";
				when "10010000111111" => data <= "000000";
				when "10010001000000" => data <= "000000";
				when "10010001000001" => data <= "000000";
				when "10010001000010" => data <= "000000";
				when "10010001000011" => data <= "000000";
				when "10010001000100" => data <= "000000";
				when "10010001000101" => data <= "000000";
				when "10010001000110" => data <= "000000";
				when "10010001000111" => data <= "000000";
				when "10010001001000" => data <= "000000";
				when "10010001001001" => data <= "000000";
				when "10010001001010" => data <= "000000";
				when "10010001001011" => data <= "000000";
				when "10010001001100" => data <= "000000";
				when "10010001001101" => data <= "000000";
				when "10010001001110" => data <= "000000";
				when "10010001001111" => data <= "000000";
				when "10010001010000" => data <= "000000";
				when "10010001010001" => data <= "000000";
				when "10010001010010" => data <= "000000";
				when "10010001010011" => data <= "000000";
				when "10010001010100" => data <= "000000";
				when "10010001010101" => data <= "000000";
				when "10010001010110" => data <= "000000";
				when "10010001010111" => data <= "000000";
				when "10010001011000" => data <= "000000";
				when "10010001011001" => data <= "000000";
				when "10010001011010" => data <= "000000";
				when "10010001011011" => data <= "000000";
				when "10010001011100" => data <= "000000";
				when "10010001011101" => data <= "000000";
				when "10010001011110" => data <= "000000";
				when "10010001011111" => data <= "000000";
				when "10010001100000" => data <= "000000";
				when "10010001100001" => data <= "000000";
				when "10010001100010" => data <= "000000";
				when "10010001100011" => data <= "000000";
				when "10010001100100" => data <= "000000";
				when "10010001100101" => data <= "000000";
				when "10010001100110" => data <= "000000";
				when "10010001100111" => data <= "000000";
				when "10010001101000" => data <= "000000";
				when "10010001101001" => data <= "000000";
				when "10010001101010" => data <= "000000";
				when "10010001101011" => data <= "000000";
				when "10010001101100" => data <= "000000";
				when "10010001101101" => data <= "000000";
				when "10010001101110" => data <= "000000";
				when "10010001101111" => data <= "000000";
				when "10010001110000" => data <= "000000";
				when "10010001110001" => data <= "000000";
				when "10010001110010" => data <= "000000";
				when "10010001110011" => data <= "000000";
				when "10010001110100" => data <= "000000";
				when "10010001110101" => data <= "000000";
				when "10010001110110" => data <= "000000";
				when "10010001110111" => data <= "000000";
				when "10010001111000" => data <= "000000";
				when "10010001111001" => data <= "000000";
				when "10010001111010" => data <= "000000";
				when "10010001111011" => data <= "000000";
				when "10010001111100" => data <= "000000";
				when "10010001111101" => data <= "000000";
				when "10010001111110" => data <= "000000";
				when "10010001111111" => data <= "000000";
				when "10010010000000" => data <= "000000";
				when "10010010000001" => data <= "000000";
				when "10010010000010" => data <= "000000";
				when "10010010000011" => data <= "000000";
				when "10010010000100" => data <= "000000";
				when "10010010000101" => data <= "000000";
				when "10010010000110" => data <= "000000";
				when "10010010000111" => data <= "000000";
				when "10010010001000" => data <= "000000";
				when "10010010001001" => data <= "000000";
				when "10010010001010" => data <= "000000";
				when "10010010001011" => data <= "000000";
				when "10010010001100" => data <= "000000";
				when "10010010001101" => data <= "000000";
				when "10010010001110" => data <= "000000";
				when "10010010001111" => data <= "000000";
				when "10010010010000" => data <= "000000";
				when "10010010010001" => data <= "000000";
				when "10010010010010" => data <= "000000";
				when "10010010010011" => data <= "000000";
				when "10010010010100" => data <= "000000";
				when "10010010010101" => data <= "000000";
				when "10010010010110" => data <= "000000";
				when "10010010010111" => data <= "000000";
				when "10010010011000" => data <= "000000";
				when "10010010011001" => data <= "000000";
				when "10010010011010" => data <= "000000";
				when "10010010011011" => data <= "000000";
				when "10010010011100" => data <= "000000";
				when "10010010011101" => data <= "000000";
				when "10010010011110" => data <= "000000";
				when "10010010011111" => data <= "000000";
				when "10010010100000" => data <= "000000";
				when "10010010100001" => data <= "000000";
				when "10010010100010" => data <= "000000";
				when "10010010100011" => data <= "000000";
				when "10010010100100" => data <= "000000";
				when "10010010100101" => data <= "000000";
				when "10010010100110" => data <= "000000";
				when "10010010100111" => data <= "000000";
				when "10010010101000" => data <= "000000";
				when "10010010101001" => data <= "000000";
				when "10010010101010" => data <= "000000";
				when "10010010101011" => data <= "000000";
				when "10010010101100" => data <= "000000";
				when "10010010101101" => data <= "000000";
				when "10010010101110" => data <= "000000";
				when "10010010101111" => data <= "000000";
				when "10010010110000" => data <= "000000";
				when "10010010110001" => data <= "000000";
				when "10010010110010" => data <= "000000";
				when "10010010110011" => data <= "000000";
				when "10010010110100" => data <= "000000";
				when "10010010110101" => data <= "000000";
				when "10010010110110" => data <= "000000";
				when "10010010110111" => data <= "000000";
				when "10010010111000" => data <= "000000";
				when "10010010111001" => data <= "000000";
				when "10010010111010" => data <= "000000";
				when "10010010111011" => data <= "000000";
				when "10010010111100" => data <= "000000";
				when "10010010111101" => data <= "000000";
				when "10010010111110" => data <= "000000";
				when "10010010111111" => data <= "000000";
				when "10010011000000" => data <= "000000";
				when "10010011000001" => data <= "000000";
				when "10010011000010" => data <= "000000";
				when "10010011000011" => data <= "000000";
				when "10010011000100" => data <= "000000";
				when "10010011000101" => data <= "000000";
				when "10010011000110" => data <= "000000";
				when "10010011000111" => data <= "000000";
				when "10010011001000" => data <= "000000";
				when "10010011001001" => data <= "000000";
				when "10010011001010" => data <= "000000";
				when "10010011001011" => data <= "000000";
				when "10010011001100" => data <= "000000";
				when "10010011001101" => data <= "000000";
				when "10010011001110" => data <= "000000";
				when "10010011001111" => data <= "000000";
				when "10010011010000" => data <= "000000";
				when "10010011010001" => data <= "000000";
				when "10010011010010" => data <= "000000";
				when "10010011010011" => data <= "000000";
				when "10010011010100" => data <= "000000";
				when "10010011010101" => data <= "000000";
				when "10010011010110" => data <= "000000";
				when "10010011010111" => data <= "000000";
				when "10010011011000" => data <= "000000";
				when "10010011011001" => data <= "000000";
				when "10010011011010" => data <= "000000";
				when "10010011011011" => data <= "000000";
				when "10010011011100" => data <= "000000";
				when "10010011011101" => data <= "000000";
				when "10010011011110" => data <= "000000";
				when "10010011011111" => data <= "000000";
				when "10010011100000" => data <= "000000";
				when "10010011100001" => data <= "000000";
				when "10010011100010" => data <= "000000";
				when "10010011100011" => data <= "000000";
				when "10010011100100" => data <= "000000";
				when "10010011100101" => data <= "000000";
				when "10010011100110" => data <= "000000";
				when "10010011100111" => data <= "000000";
				when "10010011101000" => data <= "000000";
				when "10010011101001" => data <= "000000";
				when "10010011101010" => data <= "000000";
				when "10010011101011" => data <= "000000";
				when "10010011101100" => data <= "000000";
				when "10010011101101" => data <= "000000";
				when "10010011101110" => data <= "000000";
				when "10010011101111" => data <= "000000";
				when "10010011110000" => data <= "000000";
				when "10010011110001" => data <= "000000";
				when "10010011110010" => data <= "000000";
				when "10010011110011" => data <= "000000";
				when "10010011110100" => data <= "000000";
				when "10010011110101" => data <= "000000";
				when "10010011110110" => data <= "000000";
				when "10010011110111" => data <= "000000";
				when "10010011111000" => data <= "000000";
				when "10010011111001" => data <= "000000";
				when "10010011111010" => data <= "000000";
				when "10010011111011" => data <= "000000";
				when "10010011111100" => data <= "000000";
				when "10010011111101" => data <= "000000";
				when "10010011111110" => data <= "000000";
				when "10010011111111" => data <= "000000";
				when "10010100000000" => data <= "000000";
				when "10010100000001" => data <= "000000";
				when "10010100000010" => data <= "000000";
				when "10010100000011" => data <= "000000";
				when "10010100000100" => data <= "000000";
				when "10010100000101" => data <= "000000";
				when "10010100000110" => data <= "000000";
				when "10010100000111" => data <= "000000";
				when "10010100001000" => data <= "000000";
				when "10010100001001" => data <= "000000";
				when "10010100001010" => data <= "000000";
				when "10010100001011" => data <= "000000";
				when "10010100001100" => data <= "000000";
				when "10010100001101" => data <= "000000";
				when "10010100001110" => data <= "000000";
				when "10010100001111" => data <= "000000";
				when "10010100010000" => data <= "000000";
				when "10010100010001" => data <= "000000";
				when "10010100010010" => data <= "000000";
				when "10010100010011" => data <= "000000";
				when "10010100010100" => data <= "000000";
				when "10010100010101" => data <= "000000";
				when "10010100010110" => data <= "000000";
				when "10010100010111" => data <= "000000";
				when "10010100011000" => data <= "000000";
				when "10010100011001" => data <= "000000";
				when "10010100011010" => data <= "000000";
				when "10010100011011" => data <= "000000";
				when "10010100011100" => data <= "000000";
				when "10010100011101" => data <= "000000";
				when "10010100011110" => data <= "000000";
				when "10010100011111" => data <= "000000";
				when "10010100100000" => data <= "000000";
				when "10010100100001" => data <= "000000";
				when "10010100100010" => data <= "000000";
				when "10010100100011" => data <= "000000";
				when "10010100100100" => data <= "000000";
				when "10010100100101" => data <= "000000";
				when "10010100100110" => data <= "000000";
				when "10010100100111" => data <= "000000";
				when "10010100101000" => data <= "000000";
				when "10010100101001" => data <= "000000";
				when "10010100101010" => data <= "000000";
				when "10010100101011" => data <= "000000";
				when "10010100101100" => data <= "000000";
				when "10010100101101" => data <= "000000";
				when "10010100101110" => data <= "000000";
				when "10010100101111" => data <= "000000";
				when "10010100110000" => data <= "000000";
				when "10010100110001" => data <= "000000";
				when "10010100110010" => data <= "000000";
				when "10010100110011" => data <= "000000";
				when "10010100110100" => data <= "000000";
				when "10010100110101" => data <= "000000";
				when "10010100110110" => data <= "000000";
				when "10010100110111" => data <= "000000";
				when "10010100111000" => data <= "000000";
				when "10010100111001" => data <= "000000";
				when "10010100111010" => data <= "000000";
				when "10010100111011" => data <= "000000";
				when "10010100111100" => data <= "000000";
				when "10010100111101" => data <= "000000";
				when "10010100111110" => data <= "000000";
				when "10010100111111" => data <= "000000";
				when "10010101000000" => data <= "000000";
				when "10010101000001" => data <= "000000";
				when "10010101000010" => data <= "000000";
				when "10010101000011" => data <= "000000";
				when "10010101000100" => data <= "000000";
				when "10010101000101" => data <= "000000";
				when "10010101000110" => data <= "000000";
				when "10010101000111" => data <= "000000";
				when "10010101001000" => data <= "000000";
				when "10010101001001" => data <= "000000";
				when "10010101001010" => data <= "000000";
				when "10010101001011" => data <= "000000";
				when "10010101001100" => data <= "000000";
				when "10010101001101" => data <= "000000";
				when "10010101001110" => data <= "000000";
				when "10010101001111" => data <= "000000";
				when "10010101010000" => data <= "000000";
				when "10010101010001" => data <= "000000";
				when "10010101010010" => data <= "000000";
				when "10010101010011" => data <= "000000";
				when "10010101010100" => data <= "000000";
				when "10010101010101" => data <= "000000";
				when "10010101010110" => data <= "000000";
				when "10010101010111" => data <= "000000";
				when "10010101011000" => data <= "000000";
				when "10010101011001" => data <= "000000";
				when "10010101011010" => data <= "000000";
				when "10010101011011" => data <= "000000";
				when "10010101011100" => data <= "000000";
				when "10010101011101" => data <= "000000";
				when "10010101011110" => data <= "000000";
				when "10010101011111" => data <= "000000";
				when "10010101100000" => data <= "000000";
				when "10010101100001" => data <= "000000";
				when "10010101100010" => data <= "000000";
				when "10010101100011" => data <= "000000";
				when "10010101100100" => data <= "000000";
				when "10010101100101" => data <= "000000";
				when "10010101100110" => data <= "000000";
				when "10010101100111" => data <= "000000";
				when "10010101101000" => data <= "000000";
				when "10010101101001" => data <= "000000";
				when "10010101101010" => data <= "000000";
				when "10010101101011" => data <= "000000";
				when "10010101101100" => data <= "000000";
				when "10010101101101" => data <= "000000";
				when "10010101101110" => data <= "000000";
				when "10010101101111" => data <= "000000";
				when "10010101110000" => data <= "000000";
				when "10010101110001" => data <= "000000";
				when "10010101110010" => data <= "000000";
				when "10010101110011" => data <= "000000";
				when "10010101110100" => data <= "000000";
				when "10010101110101" => data <= "000000";
				when "10010101110110" => data <= "000000";
				when "10010101110111" => data <= "000000";
				when "10010101111000" => data <= "000000";
				when "10010101111001" => data <= "000000";
				when "10010101111010" => data <= "000000";
				when "10010101111011" => data <= "000000";
				when "10010101111100" => data <= "000000";
				when "10010101111101" => data <= "000000";
				when "10010101111110" => data <= "000000";
				when "10010101111111" => data <= "000000";
				when "10010110000000" => data <= "000000";
				when "10010110000001" => data <= "000000";
				when "10010110000010" => data <= "000000";
				when "10010110000011" => data <= "000000";
				when "10010110000100" => data <= "000000";
				when "10010110000101" => data <= "000000";
				when "10010110000110" => data <= "000000";
				when "10010110000111" => data <= "000000";
				when "10010110001000" => data <= "000000";
				when "10010110001001" => data <= "000000";
				when "10010110001010" => data <= "000000";
				when "10010110001011" => data <= "000000";
				when "10010110001100" => data <= "000000";
				when "10010110001101" => data <= "000000";
				when "10010110001110" => data <= "000000";
				when "10010110001111" => data <= "000000";
				when "10010110010000" => data <= "000000";
				when "10010110010001" => data <= "000000";
				when "10010110010010" => data <= "000000";
				when "10010110010011" => data <= "000000";
				when "10010110010100" => data <= "000000";
				when "10010110010101" => data <= "000000";
				when "10010110010110" => data <= "000000";
				when "10010110010111" => data <= "000000";
				when "10010110011000" => data <= "000000";
				when "10010110011001" => data <= "000000";
				when "10010110011010" => data <= "000000";
				when "10010110011011" => data <= "000000";
				when "10010110011100" => data <= "000000";
				when "10010110011101" => data <= "000000";
				when "10010110011110" => data <= "000000";
				when "10010110011111" => data <= "000000";
				when "10010110100000" => data <= "000000";
				when "10010110100001" => data <= "000000";
				when "10010110100010" => data <= "000000";
				when "10010110100011" => data <= "000000";
				when "10010110100100" => data <= "000000";
				when "10010110100101" => data <= "000000";
				when "10010110100110" => data <= "000000";
				when "10010110100111" => data <= "000000";
				when "10010110101000" => data <= "000000";
				when "10010110101001" => data <= "000000";
				when "10010110101010" => data <= "000000";
				when "10010110101011" => data <= "000000";
				when "10010110101100" => data <= "000000";
				when "10010110101101" => data <= "000000";
				when "10010110101110" => data <= "000000";
				when "10010110101111" => data <= "000000";
				when "10010110110000" => data <= "000000";
				when "10010110110001" => data <= "000000";
				when "10010110110010" => data <= "000000";
				when "10010110110011" => data <= "000000";
				when "10010110110100" => data <= "000000";
				when "10010110110101" => data <= "000000";
				when "10010110110110" => data <= "000000";
				when "10010110110111" => data <= "000000";
				when "10010110111000" => data <= "000000";
				when "10010110111001" => data <= "000000";
				when "10010110111010" => data <= "000000";
				when "10010110111011" => data <= "000000";
				when "10010110111100" => data <= "000000";
				when "10010110111101" => data <= "000000";
				when "10010110111110" => data <= "000000";
				when "10010110111111" => data <= "000000";
				when "10010111000000" => data <= "000000";
				when "10010111000001" => data <= "000000";
				when "10010111000010" => data <= "000000";
				when "10010111000011" => data <= "000000";
				when "10010111000100" => data <= "000000";
				when "10010111000101" => data <= "000000";
				when "10010111000110" => data <= "000000";
				when "10010111000111" => data <= "000000";
				when "10010111001000" => data <= "000000";
				when "10010111001001" => data <= "000000";
				when "10010111001010" => data <= "000000";
				when "10010111001011" => data <= "000000";
				when "10010111001100" => data <= "000000";
				when "10010111001101" => data <= "000000";
				when "10010111001110" => data <= "000000";
				when "10010111001111" => data <= "000000";
				when "10010111010000" => data <= "000000";
				when "10010111010001" => data <= "000000";
				when "10010111010010" => data <= "000000";
				when "10010111010011" => data <= "000000";
				when "10010111010100" => data <= "000000";
				when "10010111010101" => data <= "000000";
				when "10010111010110" => data <= "000000";
				when "10010111010111" => data <= "000000";
				when "10010111011000" => data <= "000000";
				when "10010111011001" => data <= "000000";
				when "10010111011010" => data <= "000000";
				when "10010111011011" => data <= "000000";
				when "10010111011100" => data <= "000000";
				when "10010111011101" => data <= "000000";
				when "10010111011110" => data <= "000000";
				when "10010111011111" => data <= "000000";
				when "10010111100000" => data <= "000000";
				when "10010111100001" => data <= "000000";
				when "10010111100010" => data <= "000000";
				when "10010111100011" => data <= "000000";
				when "10010111100100" => data <= "000000";
				when "10010111100101" => data <= "000000";
				when "10010111100110" => data <= "000000";
				when "10010111100111" => data <= "000000";
				when "10010111101000" => data <= "000000";
				when "10010111101001" => data <= "000000";
				when "10010111101010" => data <= "000000";
				when "10010111101011" => data <= "000000";
				when "10010111101100" => data <= "000000";
				when "10010111101101" => data <= "000000";
				when "10010111101110" => data <= "000000";
				when "10010111101111" => data <= "000000";
				when "10010111110000" => data <= "000000";
				when "10010111110001" => data <= "000000";
				when "10010111110010" => data <= "000000";
				when "10010111110011" => data <= "000000";
				when "10010111110100" => data <= "000000";
				when "10010111110101" => data <= "000000";
				when "10010111110110" => data <= "000000";
				when "10010111110111" => data <= "000000";
				when "10010111111000" => data <= "000000";
				when "10010111111001" => data <= "000000";
				when "10010111111010" => data <= "000000";
				when "10010111111011" => data <= "000000";
				when "10010111111100" => data <= "000000";
				when "10010111111101" => data <= "000000";
				when "10010111111110" => data <= "000000";
				when "10010111111111" => data <= "000000";
				when "10011000000000" => data <= "000000";
				when "10011000000001" => data <= "000000";
				when "10011000000010" => data <= "000000";
				when "10011000000011" => data <= "000000";
				when "10011000000100" => data <= "000000";
				when "10011000000101" => data <= "000000";
				when "10011000000110" => data <= "000000";
				when "10011000000111" => data <= "000000";
				when "10011000001000" => data <= "000000";
				when "10011000001001" => data <= "000000";
				when "10011000001010" => data <= "000000";
				when "10011000001011" => data <= "000000";
				when "10011000001100" => data <= "000000";
				when "10011000001101" => data <= "000000";
				when "10011000001110" => data <= "111111";
				when "10011000001111" => data <= "111111";
				when "10011000010000" => data <= "111111";
				when "10011000010001" => data <= "111111";
				when "10011000010010" => data <= "111111";
				when "10011000010011" => data <= "000000";
				when "10011000010100" => data <= "000000";
				when "10011000010101" => data <= "000000";
				when "10011000010110" => data <= "000000";
				when "10011000010111" => data <= "111111";
				when "10011000011000" => data <= "111111";
				when "10011000011001" => data <= "111111";
				when "10011000011010" => data <= "111111";
				when "10011000011011" => data <= "111111";
				when "10011000011100" => data <= "111111";
				when "10011000011101" => data <= "000000";
				when "10011000011110" => data <= "000000";
				when "10011000011111" => data <= "000000";
				when "10011000100000" => data <= "111111";
				when "10011000100001" => data <= "111111";
				when "10011000100010" => data <= "111111";
				when "10011000100011" => data <= "111111";
				when "10011000100100" => data <= "111111";
				when "10011000100101" => data <= "111111";
				when "10011000100110" => data <= "111111";
				when "10011000100111" => data <= "000000";
				when "10011000101000" => data <= "000000";
				when "10011000101001" => data <= "000000";
				when "10011000101010" => data <= "111111";
				when "10011000101011" => data <= "111111";
				when "10011000101100" => data <= "111111";
				when "10011000101101" => data <= "111111";
				when "10011000101110" => data <= "111111";
				when "10011000101111" => data <= "111111";
				when "10011000110000" => data <= "000000";
				when "10011000110001" => data <= "000000";
				when "10011000110010" => data <= "000000";
				when "10011000110011" => data <= "000000";
				when "10011000110100" => data <= "111111";
				when "10011000110101" => data <= "111111";
				when "10011000110110" => data <= "111111";
				when "10011000110111" => data <= "111111";
				when "10011000111000" => data <= "111111";
				when "10011000111001" => data <= "111111";
				when "10011000111010" => data <= "111111";
				when "10011000111011" => data <= "000000";
				when "10011000111100" => data <= "000000";
				when "10011000111101" => data <= "000000";
				when "10011000111110" => data <= "000000";
				when "10011000111111" => data <= "000000";
				when "10011001000000" => data <= "000000";
				when "10011001000001" => data <= "000000";
				when "10011001000010" => data <= "000000";
				when "10011001000011" => data <= "000000";
				when "10011001000100" => data <= "000000";
				when "10011001000101" => data <= "111111";
				when "10011001000110" => data <= "111111";
				when "10011001000111" => data <= "111111";
				when "10011001001000" => data <= "111111";
				when "10011001001001" => data <= "111111";
				when "10011001001010" => data <= "111111";
				when "10011001001011" => data <= "111111";
				when "10011001001100" => data <= "000000";
				when "10011001001101" => data <= "000000";
				when "10011001001110" => data <= "111111";
				when "10011001001111" => data <= "111111";
				when "10011001010000" => data <= "111111";
				when "10011001010001" => data <= "111111";
				when "10011001010010" => data <= "111111";
				when "10011001010011" => data <= "111111";
				when "10011001010100" => data <= "111111";
				when "10011001010101" => data <= "111111";
				when "10011001010110" => data <= "000000";
				when "10011001010111" => data <= "000000";
				when "10011001011000" => data <= "000000";
				when "10011001011001" => data <= "000000";
				when "10011001011010" => data <= "111111";
				when "10011001011011" => data <= "111111";
				when "10011001011100" => data <= "000000";
				when "10011001011101" => data <= "000000";
				when "10011001011110" => data <= "000000";
				when "10011001011111" => data <= "000000";
				when "10011001100000" => data <= "000000";
				when "10011001100001" => data <= "000000";
				when "10011001100010" => data <= "000000";
				when "10011001100011" => data <= "000000";
				when "10011001100100" => data <= "111111";
				when "10011001100101" => data <= "111111";
				when "10011001100110" => data <= "111111";
				when "10011001100111" => data <= "111111";
				when "10011001101000" => data <= "111111";
				when "10011001101001" => data <= "111111";
				when "10011001101010" => data <= "000000";
				when "10011001101011" => data <= "000000";
				when "10011001101100" => data <= "000000";
				when "10011001101101" => data <= "111111";
				when "10011001101110" => data <= "111111";
				when "10011001101111" => data <= "111111";
				when "10011001110000" => data <= "111111";
				when "10011001110001" => data <= "111111";
				when "10011001110010" => data <= "111111";
				when "10011001110011" => data <= "111111";
				when "10011001110100" => data <= "111111";
				when "10011001110101" => data <= "000000";
				when "10011001110110" => data <= "000000";
				when "10011001110111" => data <= "000000";
				when "10011001111000" => data <= "000000";
				when "10011001111001" => data <= "000000";
				when "10011001111010" => data <= "000000";
				when "10011001111011" => data <= "000000";
				when "10011001111100" => data <= "000000";
				when "10011001111101" => data <= "000000";
				when "10011001111110" => data <= "000000";
				when "10011001111111" => data <= "000000";
				when "10011010000000" => data <= "000000";
				when "10011010000001" => data <= "000000";
				when "10011010000010" => data <= "000000";
				when "10011010000011" => data <= "000000";
				when "10011010000100" => data <= "000000";
				when "10011010000101" => data <= "000000";
				when "10011010000110" => data <= "000000";
				when "10011010000111" => data <= "000000";
				when "10011010001000" => data <= "000000";
				when "10011010001001" => data <= "000000";
				when "10011010001010" => data <= "000000";
				when "10011010001011" => data <= "000000";
				when "10011010001100" => data <= "000000";
				when "10011010001101" => data <= "111111";
				when "10011010001110" => data <= "111111";
				when "10011010001111" => data <= "111111";
				when "10011010010000" => data <= "111111";
				when "10011010010001" => data <= "111111";
				when "10011010010010" => data <= "111111";
				when "10011010010011" => data <= "000000";
				when "10011010010100" => data <= "000000";
				when "10011010010101" => data <= "000000";
				when "10011010010110" => data <= "111111";
				when "10011010010111" => data <= "111111";
				when "10011010011000" => data <= "111111";
				when "10011010011001" => data <= "111111";
				when "10011010011010" => data <= "111111";
				when "10011010011011" => data <= "111111";
				when "10011010011100" => data <= "111111";
				when "10011010011101" => data <= "111111";
				when "10011010011110" => data <= "000000";
				when "10011010011111" => data <= "000000";
				when "10011010100000" => data <= "111111";
				when "10011010100001" => data <= "111111";
				when "10011010100010" => data <= "111111";
				when "10011010100011" => data <= "111111";
				when "10011010100100" => data <= "111111";
				when "10011010100101" => data <= "111111";
				when "10011010100110" => data <= "111111";
				when "10011010100111" => data <= "000000";
				when "10011010101000" => data <= "000000";
				when "10011010101001" => data <= "000000";
				when "10011010101010" => data <= "111111";
				when "10011010101011" => data <= "111111";
				when "10011010101100" => data <= "111111";
				when "10011010101101" => data <= "111111";
				when "10011010101110" => data <= "111111";
				when "10011010101111" => data <= "111111";
				when "10011010110000" => data <= "000000";
				when "10011010110001" => data <= "000000";
				when "10011010110010" => data <= "000000";
				when "10011010110011" => data <= "000000";
				when "10011010110100" => data <= "111111";
				when "10011010110101" => data <= "111111";
				when "10011010110110" => data <= "111111";
				when "10011010110111" => data <= "111111";
				when "10011010111000" => data <= "111111";
				when "10011010111001" => data <= "111111";
				when "10011010111010" => data <= "111111";
				when "10011010111011" => data <= "000000";
				when "10011010111100" => data <= "000000";
				when "10011010111101" => data <= "000000";
				when "10011010111110" => data <= "000000";
				when "10011010111111" => data <= "000000";
				when "10011011000000" => data <= "000000";
				when "10011011000001" => data <= "000000";
				when "10011011000010" => data <= "000000";
				when "10011011000011" => data <= "000000";
				when "10011011000100" => data <= "000000";
				when "10011011000101" => data <= "111111";
				when "10011011000110" => data <= "111111";
				when "10011011000111" => data <= "111111";
				when "10011011001000" => data <= "111111";
				when "10011011001001" => data <= "111111";
				when "10011011001010" => data <= "111111";
				when "10011011001011" => data <= "111111";
				when "10011011001100" => data <= "000000";
				when "10011011001101" => data <= "000000";
				when "10011011001110" => data <= "111111";
				when "10011011001111" => data <= "111111";
				when "10011011010000" => data <= "111111";
				when "10011011010001" => data <= "111111";
				when "10011011010010" => data <= "111111";
				when "10011011010011" => data <= "111111";
				when "10011011010100" => data <= "111111";
				when "10011011010101" => data <= "111111";
				when "10011011010110" => data <= "000000";
				when "10011011010111" => data <= "000000";
				when "10011011011000" => data <= "000000";
				when "10011011011001" => data <= "000000";
				when "10011011011010" => data <= "111111";
				when "10011011011011" => data <= "111111";
				when "10011011011100" => data <= "000000";
				when "10011011011101" => data <= "000000";
				when "10011011011110" => data <= "000000";
				when "10011011011111" => data <= "000000";
				when "10011011100000" => data <= "000000";
				when "10011011100001" => data <= "000000";
				when "10011011100010" => data <= "000000";
				when "10011011100011" => data <= "111111";
				when "10011011100100" => data <= "111111";
				when "10011011100101" => data <= "111111";
				when "10011011100110" => data <= "111111";
				when "10011011100111" => data <= "111111";
				when "10011011101000" => data <= "111111";
				when "10011011101001" => data <= "111111";
				when "10011011101010" => data <= "111111";
				when "10011011101011" => data <= "000000";
				when "10011011101100" => data <= "000000";
				when "10011011101101" => data <= "111111";
				when "10011011101110" => data <= "111111";
				when "10011011101111" => data <= "111111";
				when "10011011110000" => data <= "111111";
				when "10011011110001" => data <= "111111";
				when "10011011110010" => data <= "111111";
				when "10011011110011" => data <= "111111";
				when "10011011110100" => data <= "111111";
				when "10011011110101" => data <= "000000";
				when "10011011110110" => data <= "000000";
				when "10011011110111" => data <= "000000";
				when "10011011111000" => data <= "000000";
				when "10011011111001" => data <= "000000";
				when "10011011111010" => data <= "000000";
				when "10011011111011" => data <= "000000";
				when "10011011111100" => data <= "000000";
				when "10011011111101" => data <= "000000";
				when "10011011111110" => data <= "000000";
				when "10011011111111" => data <= "000000";
				when "10011100000000" => data <= "000000";
				when "10011100000001" => data <= "000000";
				when "10011100000010" => data <= "000000";
				when "10011100000011" => data <= "000000";
				when "10011100000100" => data <= "000000";
				when "10011100000101" => data <= "000000";
				when "10011100000110" => data <= "000000";
				when "10011100000111" => data <= "000000";
				when "10011100001000" => data <= "000000";
				when "10011100001001" => data <= "000000";
				when "10011100001010" => data <= "000000";
				when "10011100001011" => data <= "000000";
				when "10011100001100" => data <= "000000";
				when "10011100001101" => data <= "111111";
				when "10011100001110" => data <= "111111";
				when "10011100001111" => data <= "000000";
				when "10011100010000" => data <= "000000";
				when "10011100010001" => data <= "000000";
				when "10011100010010" => data <= "000000";
				when "10011100010011" => data <= "111111";
				when "10011100010100" => data <= "111111";
				when "10011100010101" => data <= "000000";
				when "10011100010110" => data <= "111111";
				when "10011100010111" => data <= "111111";
				when "10011100011000" => data <= "000000";
				when "10011100011001" => data <= "000000";
				when "10011100011010" => data <= "000000";
				when "10011100011011" => data <= "000000";
				when "10011100011100" => data <= "111111";
				when "10011100011101" => data <= "111111";
				when "10011100011110" => data <= "000000";
				when "10011100011111" => data <= "000000";
				when "10011100100000" => data <= "111111";
				when "10011100100001" => data <= "111111";
				when "10011100100010" => data <= "000000";
				when "10011100100011" => data <= "000000";
				when "10011100100100" => data <= "000000";
				when "10011100100101" => data <= "000000";
				when "10011100100110" => data <= "000000";
				when "10011100100111" => data <= "000000";
				when "10011100101000" => data <= "111111";
				when "10011100101001" => data <= "111111";
				when "10011100101010" => data <= "000000";
				when "10011100101011" => data <= "000000";
				when "10011100101100" => data <= "000000";
				when "10011100101101" => data <= "000000";
				when "10011100101110" => data <= "000000";
				when "10011100101111" => data <= "000000";
				when "10011100110000" => data <= "000000";
				when "10011100110001" => data <= "000000";
				when "10011100110010" => data <= "111111";
				when "10011100110011" => data <= "111111";
				when "10011100110100" => data <= "000000";
				when "10011100110101" => data <= "000000";
				when "10011100110110" => data <= "000000";
				when "10011100110111" => data <= "000000";
				when "10011100111000" => data <= "000000";
				when "10011100111001" => data <= "000000";
				when "10011100111010" => data <= "000000";
				when "10011100111011" => data <= "000000";
				when "10011100111100" => data <= "000000";
				when "10011100111101" => data <= "000000";
				when "10011100111110" => data <= "000000";
				when "10011100111111" => data <= "000000";
				when "10011101000000" => data <= "000000";
				when "10011101000001" => data <= "000000";
				when "10011101000010" => data <= "000000";
				when "10011101000011" => data <= "000000";
				when "10011101000100" => data <= "111111";
				when "10011101000101" => data <= "111111";
				when "10011101000110" => data <= "000000";
				when "10011101000111" => data <= "000000";
				when "10011101001000" => data <= "000000";
				when "10011101001001" => data <= "000000";
				when "10011101001010" => data <= "000000";
				when "10011101001011" => data <= "000000";
				when "10011101001100" => data <= "000000";
				when "10011101001101" => data <= "000000";
				when "10011101001110" => data <= "000000";
				when "10011101001111" => data <= "000000";
				when "10011101010000" => data <= "000000";
				when "10011101010001" => data <= "111111";
				when "10011101010010" => data <= "111111";
				when "10011101010011" => data <= "000000";
				when "10011101010100" => data <= "000000";
				when "10011101010101" => data <= "000000";
				when "10011101010110" => data <= "000000";
				when "10011101010111" => data <= "000000";
				when "10011101011000" => data <= "111111";
				when "10011101011001" => data <= "111111";
				when "10011101011010" => data <= "000000";
				when "10011101011011" => data <= "000000";
				when "10011101011100" => data <= "111111";
				when "10011101011101" => data <= "111111";
				when "10011101011110" => data <= "000000";
				when "10011101011111" => data <= "000000";
				when "10011101100000" => data <= "000000";
				when "10011101100001" => data <= "000000";
				when "10011101100010" => data <= "000000";
				when "10011101100011" => data <= "111111";
				when "10011101100100" => data <= "111111";
				when "10011101100101" => data <= "000000";
				when "10011101100110" => data <= "000000";
				when "10011101100111" => data <= "000000";
				when "10011101101000" => data <= "000000";
				when "10011101101001" => data <= "111111";
				when "10011101101010" => data <= "111111";
				when "10011101101011" => data <= "000000";
				when "10011101101100" => data <= "000000";
				when "10011101101101" => data <= "000000";
				when "10011101101110" => data <= "000000";
				when "10011101101111" => data <= "000000";
				when "10011101110000" => data <= "111111";
				when "10011101110001" => data <= "111111";
				when "10011101110010" => data <= "000000";
				when "10011101110011" => data <= "000000";
				when "10011101110100" => data <= "000000";
				when "10011101110101" => data <= "000000";
				when "10011101110110" => data <= "000000";
				when "10011101110111" => data <= "000000";
				when "10011101111000" => data <= "000000";
				when "10011101111001" => data <= "000000";
				when "10011101111010" => data <= "000000";
				when "10011101111011" => data <= "000000";
				when "10011101111100" => data <= "000000";
				when "10011101111101" => data <= "000000";
				when "10011101111110" => data <= "000000";
				when "10011101111111" => data <= "000000";
				when "10011110000000" => data <= "000000";
				when "10011110000001" => data <= "000000";
				when "10011110000010" => data <= "000000";
				when "10011110000011" => data <= "000000";
				when "10011110000100" => data <= "000000";
				when "10011110000101" => data <= "000000";
				when "10011110000110" => data <= "000000";
				when "10011110000111" => data <= "000000";
				when "10011110001000" => data <= "000000";
				when "10011110001001" => data <= "000000";
				when "10011110001010" => data <= "000000";
				when "10011110001011" => data <= "000000";
				when "10011110001100" => data <= "000000";
				when "10011110001101" => data <= "111111";
				when "10011110001110" => data <= "111111";
				when "10011110001111" => data <= "000000";
				when "10011110010000" => data <= "000000";
				when "10011110010001" => data <= "000000";
				when "10011110010010" => data <= "000000";
				when "10011110010011" => data <= "111111";
				when "10011110010100" => data <= "111111";
				when "10011110010101" => data <= "000000";
				when "10011110010110" => data <= "111111";
				when "10011110010111" => data <= "111111";
				when "10011110011000" => data <= "000000";
				when "10011110011001" => data <= "000000";
				when "10011110011010" => data <= "000000";
				when "10011110011011" => data <= "000000";
				when "10011110011100" => data <= "111111";
				when "10011110011101" => data <= "111111";
				when "10011110011110" => data <= "000000";
				when "10011110011111" => data <= "000000";
				when "10011110100000" => data <= "111111";
				when "10011110100001" => data <= "111111";
				when "10011110100010" => data <= "000000";
				when "10011110100011" => data <= "000000";
				when "10011110100100" => data <= "000000";
				when "10011110100101" => data <= "000000";
				when "10011110100110" => data <= "000000";
				when "10011110100111" => data <= "000000";
				when "10011110101000" => data <= "111111";
				when "10011110101001" => data <= "111111";
				when "10011110101010" => data <= "000000";
				when "10011110101011" => data <= "000000";
				when "10011110101100" => data <= "000000";
				when "10011110101101" => data <= "000000";
				when "10011110101110" => data <= "000000";
				when "10011110101111" => data <= "000000";
				when "10011110110000" => data <= "000000";
				when "10011110110001" => data <= "000000";
				when "10011110110010" => data <= "111111";
				when "10011110110011" => data <= "111111";
				when "10011110110100" => data <= "000000";
				when "10011110110101" => data <= "000000";
				when "10011110110110" => data <= "000000";
				when "10011110110111" => data <= "000000";
				when "10011110111000" => data <= "000000";
				when "10011110111001" => data <= "000000";
				when "10011110111010" => data <= "000000";
				when "10011110111011" => data <= "000000";
				when "10011110111100" => data <= "000000";
				when "10011110111101" => data <= "000000";
				when "10011110111110" => data <= "000000";
				when "10011110111111" => data <= "000000";
				when "10011111000000" => data <= "000000";
				when "10011111000001" => data <= "000000";
				when "10011111000010" => data <= "000000";
				when "10011111000011" => data <= "000000";
				when "10011111000100" => data <= "111111";
				when "10011111000101" => data <= "111111";
				when "10011111000110" => data <= "000000";
				when "10011111000111" => data <= "000000";
				when "10011111001000" => data <= "000000";
				when "10011111001001" => data <= "000000";
				when "10011111001010" => data <= "000000";
				when "10011111001011" => data <= "000000";
				when "10011111001100" => data <= "000000";
				when "10011111001101" => data <= "000000";
				when "10011111001110" => data <= "000000";
				when "10011111001111" => data <= "000000";
				when "10011111010000" => data <= "000000";
				when "10011111010001" => data <= "111111";
				when "10011111010010" => data <= "111111";
				when "10011111010011" => data <= "000000";
				when "10011111010100" => data <= "000000";
				when "10011111010101" => data <= "000000";
				when "10011111010110" => data <= "000000";
				when "10011111010111" => data <= "000000";
				when "10011111011000" => data <= "111111";
				when "10011111011001" => data <= "111111";
				when "10011111011010" => data <= "000000";
				when "10011111011011" => data <= "000000";
				when "10011111011100" => data <= "111111";
				when "10011111011101" => data <= "111111";
				when "10011111011110" => data <= "000000";
				when "10011111011111" => data <= "000000";
				when "10011111100000" => data <= "000000";
				when "10011111100001" => data <= "000000";
				when "10011111100010" => data <= "000000";
				when "10011111100011" => data <= "111111";
				when "10011111100100" => data <= "111111";
				when "10011111100101" => data <= "000000";
				when "10011111100110" => data <= "000000";
				when "10011111100111" => data <= "000000";
				when "10011111101000" => data <= "000000";
				when "10011111101001" => data <= "111111";
				when "10011111101010" => data <= "111111";
				when "10011111101011" => data <= "000000";
				when "10011111101100" => data <= "000000";
				when "10011111101101" => data <= "000000";
				when "10011111101110" => data <= "000000";
				when "10011111101111" => data <= "000000";
				when "10011111110000" => data <= "111111";
				when "10011111110001" => data <= "111111";
				when "10011111110010" => data <= "000000";
				when "10011111110011" => data <= "000000";
				when "10011111110100" => data <= "000000";
				when "10011111110101" => data <= "000000";
				when "10011111110110" => data <= "000000";
				when "10011111110111" => data <= "000000";
				when "10011111111000" => data <= "000000";
				when "10011111111001" => data <= "000000";
				when "10011111111010" => data <= "000000";
				when "10011111111011" => data <= "000000";
				when "10011111111100" => data <= "000000";
				when "10011111111101" => data <= "000000";
				when "10011111111110" => data <= "000000";
				when "10011111111111" => data <= "000000";
				when "10100000000000" => data <= "000000";
				when "10100000000001" => data <= "000000";
				when "10100000000010" => data <= "000000";
				when "10100000000011" => data <= "000000";
				when "10100000000100" => data <= "000000";
				when "10100000000101" => data <= "000000";
				when "10100000000110" => data <= "000000";
				when "10100000000111" => data <= "000000";
				when "10100000001000" => data <= "000000";
				when "10100000001001" => data <= "000000";
				when "10100000001010" => data <= "000000";
				when "10100000001011" => data <= "000000";
				when "10100000001100" => data <= "000000";
				when "10100000001101" => data <= "111111";
				when "10100000001110" => data <= "111111";
				when "10100000001111" => data <= "000000";
				when "10100000010000" => data <= "000000";
				when "10100000010001" => data <= "000000";
				when "10100000010010" => data <= "000000";
				when "10100000010011" => data <= "111111";
				when "10100000010100" => data <= "111111";
				when "10100000010101" => data <= "000000";
				when "10100000010110" => data <= "111111";
				when "10100000010111" => data <= "111111";
				when "10100000011000" => data <= "000000";
				when "10100000011001" => data <= "000000";
				when "10100000011010" => data <= "000000";
				when "10100000011011" => data <= "000000";
				when "10100000011100" => data <= "111111";
				when "10100000011101" => data <= "111111";
				when "10100000011110" => data <= "000000";
				when "10100000011111" => data <= "000000";
				when "10100000100000" => data <= "111111";
				when "10100000100001" => data <= "111111";
				when "10100000100010" => data <= "000000";
				when "10100000100011" => data <= "000000";
				when "10100000100100" => data <= "000000";
				when "10100000100101" => data <= "000000";
				when "10100000100110" => data <= "000000";
				when "10100000100111" => data <= "000000";
				when "10100000101000" => data <= "111111";
				when "10100000101001" => data <= "111111";
				when "10100000101010" => data <= "000000";
				when "10100000101011" => data <= "000000";
				when "10100000101100" => data <= "000000";
				when "10100000101101" => data <= "000000";
				when "10100000101110" => data <= "000000";
				when "10100000101111" => data <= "000000";
				when "10100000110000" => data <= "000000";
				when "10100000110001" => data <= "000000";
				when "10100000110010" => data <= "111111";
				when "10100000110011" => data <= "111111";
				when "10100000110100" => data <= "000000";
				when "10100000110101" => data <= "000000";
				when "10100000110110" => data <= "000000";
				when "10100000110111" => data <= "000000";
				when "10100000111000" => data <= "000000";
				when "10100000111001" => data <= "000000";
				when "10100000111010" => data <= "000000";
				when "10100000111011" => data <= "000000";
				when "10100000111100" => data <= "000000";
				when "10100000111101" => data <= "000000";
				when "10100000111110" => data <= "000000";
				when "10100000111111" => data <= "000000";
				when "10100001000000" => data <= "000000";
				when "10100001000001" => data <= "000000";
				when "10100001000010" => data <= "000000";
				when "10100001000011" => data <= "000000";
				when "10100001000100" => data <= "111111";
				when "10100001000101" => data <= "111111";
				when "10100001000110" => data <= "000000";
				when "10100001000111" => data <= "000000";
				when "10100001001000" => data <= "000000";
				when "10100001001001" => data <= "000000";
				when "10100001001010" => data <= "000000";
				when "10100001001011" => data <= "000000";
				when "10100001001100" => data <= "000000";
				when "10100001001101" => data <= "000000";
				when "10100001001110" => data <= "000000";
				when "10100001001111" => data <= "000000";
				when "10100001010000" => data <= "000000";
				when "10100001010001" => data <= "111111";
				when "10100001010010" => data <= "111111";
				when "10100001010011" => data <= "000000";
				when "10100001010100" => data <= "000000";
				when "10100001010101" => data <= "000000";
				when "10100001010110" => data <= "111111";
				when "10100001010111" => data <= "111111";
				when "10100001011000" => data <= "000000";
				when "10100001011001" => data <= "000000";
				when "10100001011010" => data <= "000000";
				when "10100001011011" => data <= "000000";
				when "10100001011100" => data <= "000000";
				when "10100001011101" => data <= "000000";
				when "10100001011110" => data <= "111111";
				when "10100001011111" => data <= "111111";
				when "10100001100000" => data <= "000000";
				when "10100001100001" => data <= "000000";
				when "10100001100010" => data <= "000000";
				when "10100001100011" => data <= "111111";
				when "10100001100100" => data <= "111111";
				when "10100001100101" => data <= "000000";
				when "10100001100110" => data <= "000000";
				when "10100001100111" => data <= "000000";
				when "10100001101000" => data <= "000000";
				when "10100001101001" => data <= "111111";
				when "10100001101010" => data <= "111111";
				when "10100001101011" => data <= "000000";
				when "10100001101100" => data <= "000000";
				when "10100001101101" => data <= "000000";
				when "10100001101110" => data <= "000000";
				when "10100001101111" => data <= "000000";
				when "10100001110000" => data <= "111111";
				when "10100001110001" => data <= "111111";
				when "10100001110010" => data <= "000000";
				when "10100001110011" => data <= "000000";
				when "10100001110100" => data <= "000000";
				when "10100001110101" => data <= "000000";
				when "10100001110110" => data <= "000000";
				when "10100001110111" => data <= "000000";
				when "10100001111000" => data <= "000000";
				when "10100001111001" => data <= "000000";
				when "10100001111010" => data <= "000000";
				when "10100001111011" => data <= "000000";
				when "10100001111100" => data <= "000000";
				when "10100001111101" => data <= "000000";
				when "10100001111110" => data <= "000000";
				when "10100001111111" => data <= "000000";
				when "10100010000000" => data <= "000000";
				when "10100010000001" => data <= "000000";
				when "10100010000010" => data <= "000000";
				when "10100010000011" => data <= "000000";
				when "10100010000100" => data <= "000000";
				when "10100010000101" => data <= "000000";
				when "10100010000110" => data <= "000000";
				when "10100010000111" => data <= "000000";
				when "10100010001000" => data <= "000000";
				when "10100010001001" => data <= "000000";
				when "10100010001010" => data <= "000000";
				when "10100010001011" => data <= "000000";
				when "10100010001100" => data <= "000000";
				when "10100010001101" => data <= "111111";
				when "10100010001110" => data <= "111111";
				when "10100010001111" => data <= "000000";
				when "10100010010000" => data <= "000000";
				when "10100010010001" => data <= "000000";
				when "10100010010010" => data <= "000000";
				when "10100010010011" => data <= "111111";
				when "10100010010100" => data <= "111111";
				when "10100010010101" => data <= "000000";
				when "10100010010110" => data <= "111111";
				when "10100010010111" => data <= "111111";
				when "10100010011000" => data <= "000000";
				when "10100010011001" => data <= "000000";
				when "10100010011010" => data <= "000000";
				when "10100010011011" => data <= "000000";
				when "10100010011100" => data <= "111111";
				when "10100010011101" => data <= "111111";
				when "10100010011110" => data <= "000000";
				when "10100010011111" => data <= "000000";
				when "10100010100000" => data <= "111111";
				when "10100010100001" => data <= "111111";
				when "10100010100010" => data <= "000000";
				when "10100010100011" => data <= "000000";
				when "10100010100100" => data <= "000000";
				when "10100010100101" => data <= "000000";
				when "10100010100110" => data <= "000000";
				when "10100010100111" => data <= "000000";
				when "10100010101000" => data <= "111111";
				when "10100010101001" => data <= "111111";
				when "10100010101010" => data <= "000000";
				when "10100010101011" => data <= "000000";
				when "10100010101100" => data <= "000000";
				when "10100010101101" => data <= "000000";
				when "10100010101110" => data <= "000000";
				when "10100010101111" => data <= "000000";
				when "10100010110000" => data <= "000000";
				when "10100010110001" => data <= "000000";
				when "10100010110010" => data <= "111111";
				when "10100010110011" => data <= "111111";
				when "10100010110100" => data <= "000000";
				when "10100010110101" => data <= "000000";
				when "10100010110110" => data <= "000000";
				when "10100010110111" => data <= "000000";
				when "10100010111000" => data <= "000000";
				when "10100010111001" => data <= "000000";
				when "10100010111010" => data <= "000000";
				when "10100010111011" => data <= "000000";
				when "10100010111100" => data <= "000000";
				when "10100010111101" => data <= "000000";
				when "10100010111110" => data <= "000000";
				when "10100010111111" => data <= "000000";
				when "10100011000000" => data <= "000000";
				when "10100011000001" => data <= "000000";
				when "10100011000010" => data <= "000000";
				when "10100011000011" => data <= "000000";
				when "10100011000100" => data <= "111111";
				when "10100011000101" => data <= "111111";
				when "10100011000110" => data <= "000000";
				when "10100011000111" => data <= "000000";
				when "10100011001000" => data <= "000000";
				when "10100011001001" => data <= "000000";
				when "10100011001010" => data <= "000000";
				when "10100011001011" => data <= "000000";
				when "10100011001100" => data <= "000000";
				when "10100011001101" => data <= "000000";
				when "10100011001110" => data <= "000000";
				when "10100011001111" => data <= "000000";
				when "10100011010000" => data <= "000000";
				when "10100011010001" => data <= "111111";
				when "10100011010010" => data <= "111111";
				when "10100011010011" => data <= "000000";
				when "10100011010100" => data <= "000000";
				when "10100011010101" => data <= "000000";
				when "10100011010110" => data <= "111111";
				when "10100011010111" => data <= "111111";
				when "10100011011000" => data <= "000000";
				when "10100011011001" => data <= "000000";
				when "10100011011010" => data <= "000000";
				when "10100011011011" => data <= "000000";
				when "10100011011100" => data <= "000000";
				when "10100011011101" => data <= "000000";
				when "10100011011110" => data <= "111111";
				when "10100011011111" => data <= "111111";
				when "10100011100000" => data <= "000000";
				when "10100011100001" => data <= "000000";
				when "10100011100010" => data <= "000000";
				when "10100011100011" => data <= "111111";
				when "10100011100100" => data <= "111111";
				when "10100011100101" => data <= "000000";
				when "10100011100110" => data <= "000000";
				when "10100011100111" => data <= "000000";
				when "10100011101000" => data <= "000000";
				when "10100011101001" => data <= "111111";
				when "10100011101010" => data <= "111111";
				when "10100011101011" => data <= "000000";
				when "10100011101100" => data <= "000000";
				when "10100011101101" => data <= "000000";
				when "10100011101110" => data <= "000000";
				when "10100011101111" => data <= "000000";
				when "10100011110000" => data <= "111111";
				when "10100011110001" => data <= "111111";
				when "10100011110010" => data <= "000000";
				when "10100011110011" => data <= "000000";
				when "10100011110100" => data <= "000000";
				when "10100011110101" => data <= "000000";
				when "10100011110110" => data <= "000000";
				when "10100011110111" => data <= "000000";
				when "10100011111000" => data <= "000000";
				when "10100011111001" => data <= "000000";
				when "10100011111010" => data <= "000000";
				when "10100011111011" => data <= "000000";
				when "10100011111100" => data <= "000000";
				when "10100011111101" => data <= "000000";
				when "10100011111110" => data <= "000000";
				when "10100011111111" => data <= "000000";
				when "10100100000000" => data <= "000000";
				when "10100100000001" => data <= "000000";
				when "10100100000010" => data <= "000000";
				when "10100100000011" => data <= "000000";
				when "10100100000100" => data <= "000000";
				when "10100100000101" => data <= "000000";
				when "10100100000110" => data <= "000000";
				when "10100100000111" => data <= "000000";
				when "10100100001000" => data <= "000000";
				when "10100100001001" => data <= "000000";
				when "10100100001010" => data <= "000000";
				when "10100100001011" => data <= "000000";
				when "10100100001100" => data <= "000000";
				when "10100100001101" => data <= "111111";
				when "10100100001110" => data <= "111111";
				when "10100100001111" => data <= "111111";
				when "10100100010000" => data <= "111111";
				when "10100100010001" => data <= "111111";
				when "10100100010010" => data <= "111111";
				when "10100100010011" => data <= "000000";
				when "10100100010100" => data <= "000000";
				when "10100100010101" => data <= "000000";
				when "10100100010110" => data <= "111111";
				when "10100100010111" => data <= "111111";
				when "10100100011000" => data <= "111111";
				when "10100100011001" => data <= "111111";
				when "10100100011010" => data <= "111111";
				when "10100100011011" => data <= "111111";
				when "10100100011100" => data <= "000000";
				when "10100100011101" => data <= "000000";
				when "10100100011110" => data <= "000000";
				when "10100100011111" => data <= "000000";
				when "10100100100000" => data <= "111111";
				when "10100100100001" => data <= "111111";
				when "10100100100010" => data <= "111111";
				when "10100100100011" => data <= "111111";
				when "10100100100100" => data <= "111111";
				when "10100100100101" => data <= "000000";
				when "10100100100110" => data <= "000000";
				when "10100100100111" => data <= "000000";
				when "10100100101000" => data <= "111111";
				when "10100100101001" => data <= "111111";
				when "10100100101010" => data <= "111111";
				when "10100100101011" => data <= "111111";
				when "10100100101100" => data <= "111111";
				when "10100100101101" => data <= "111111";
				when "10100100101110" => data <= "111111";
				when "10100100101111" => data <= "111111";
				when "10100100110000" => data <= "000000";
				when "10100100110001" => data <= "000000";
				when "10100100110010" => data <= "111111";
				when "10100100110011" => data <= "111111";
				when "10100100110100" => data <= "111111";
				when "10100100110101" => data <= "111111";
				when "10100100110110" => data <= "111111";
				when "10100100110111" => data <= "111111";
				when "10100100111000" => data <= "111111";
				when "10100100111001" => data <= "111111";
				when "10100100111010" => data <= "111111";
				when "10100100111011" => data <= "000000";
				when "10100100111100" => data <= "000000";
				when "10100100111101" => data <= "000000";
				when "10100100111110" => data <= "000000";
				when "10100100111111" => data <= "000000";
				when "10100101000000" => data <= "000000";
				when "10100101000001" => data <= "000000";
				when "10100101000010" => data <= "000000";
				when "10100101000011" => data <= "000000";
				when "10100101000100" => data <= "111111";
				when "10100101000101" => data <= "111111";
				when "10100101000110" => data <= "111111";
				when "10100101000111" => data <= "111111";
				when "10100101001000" => data <= "111111";
				when "10100101001001" => data <= "111111";
				when "10100101001010" => data <= "111111";
				when "10100101001011" => data <= "111111";
				when "10100101001100" => data <= "000000";
				when "10100101001101" => data <= "000000";
				when "10100101001110" => data <= "000000";
				when "10100101001111" => data <= "000000";
				when "10100101010000" => data <= "000000";
				when "10100101010001" => data <= "111111";
				when "10100101010010" => data <= "111111";
				when "10100101010011" => data <= "000000";
				when "10100101010100" => data <= "000000";
				when "10100101010101" => data <= "000000";
				when "10100101010110" => data <= "111111";
				when "10100101010111" => data <= "111111";
				when "10100101011000" => data <= "111111";
				when "10100101011001" => data <= "111111";
				when "10100101011010" => data <= "111111";
				when "10100101011011" => data <= "111111";
				when "10100101011100" => data <= "111111";
				when "10100101011101" => data <= "111111";
				when "10100101011110" => data <= "111111";
				when "10100101011111" => data <= "111111";
				when "10100101100000" => data <= "000000";
				when "10100101100001" => data <= "000000";
				when "10100101100010" => data <= "000000";
				when "10100101100011" => data <= "111111";
				when "10100101100100" => data <= "111111";
				when "10100101100101" => data <= "111111";
				when "10100101100110" => data <= "111111";
				when "10100101100111" => data <= "111111";
				when "10100101101000" => data <= "111111";
				when "10100101101001" => data <= "000000";
				when "10100101101010" => data <= "000000";
				when "10100101101011" => data <= "000000";
				when "10100101101100" => data <= "000000";
				when "10100101101101" => data <= "000000";
				when "10100101101110" => data <= "000000";
				when "10100101101111" => data <= "000000";
				when "10100101110000" => data <= "111111";
				when "10100101110001" => data <= "111111";
				when "10100101110010" => data <= "000000";
				when "10100101110011" => data <= "000000";
				when "10100101110100" => data <= "000000";
				when "10100101110101" => data <= "000000";
				when "10100101110110" => data <= "000000";
				when "10100101110111" => data <= "000000";
				when "10100101111000" => data <= "000000";
				when "10100101111001" => data <= "000000";
				when "10100101111010" => data <= "000000";
				when "10100101111011" => data <= "000000";
				when "10100101111100" => data <= "000000";
				when "10100101111101" => data <= "000000";
				when "10100101111110" => data <= "000000";
				when "10100101111111" => data <= "000000";
				when "10100110000000" => data <= "000000";
				when "10100110000001" => data <= "000000";
				when "10100110000010" => data <= "000000";
				when "10100110000011" => data <= "000000";
				when "10100110000100" => data <= "000000";
				when "10100110000101" => data <= "000000";
				when "10100110000110" => data <= "000000";
				when "10100110000111" => data <= "000000";
				when "10100110001000" => data <= "000000";
				when "10100110001001" => data <= "000000";
				when "10100110001010" => data <= "000000";
				when "10100110001011" => data <= "000000";
				when "10100110001100" => data <= "000000";
				when "10100110001101" => data <= "111111";
				when "10100110001110" => data <= "111111";
				when "10100110001111" => data <= "111111";
				when "10100110010000" => data <= "111111";
				when "10100110010001" => data <= "111111";
				when "10100110010010" => data <= "111111";
				when "10100110010011" => data <= "000000";
				when "10100110010100" => data <= "000000";
				when "10100110010101" => data <= "000000";
				when "10100110010110" => data <= "111111";
				when "10100110010111" => data <= "111111";
				when "10100110011000" => data <= "111111";
				when "10100110011001" => data <= "111111";
				when "10100110011010" => data <= "111111";
				when "10100110011011" => data <= "111111";
				when "10100110011100" => data <= "111111";
				when "10100110011101" => data <= "111111";
				when "10100110011110" => data <= "000000";
				when "10100110011111" => data <= "000000";
				when "10100110100000" => data <= "111111";
				when "10100110100001" => data <= "111111";
				when "10100110100010" => data <= "111111";
				when "10100110100011" => data <= "111111";
				when "10100110100100" => data <= "111111";
				when "10100110100101" => data <= "000000";
				when "10100110100110" => data <= "000000";
				when "10100110100111" => data <= "000000";
				when "10100110101000" => data <= "000000";
				when "10100110101001" => data <= "000000";
				when "10100110101010" => data <= "111111";
				when "10100110101011" => data <= "111111";
				when "10100110101100" => data <= "111111";
				when "10100110101101" => data <= "111111";
				when "10100110101110" => data <= "111111";
				when "10100110101111" => data <= "111111";
				when "10100110110000" => data <= "111111";
				when "10100110110001" => data <= "000000";
				when "10100110110010" => data <= "000000";
				when "10100110110011" => data <= "000000";
				when "10100110110100" => data <= "111111";
				when "10100110110101" => data <= "111111";
				when "10100110110110" => data <= "111111";
				when "10100110110111" => data <= "111111";
				when "10100110111000" => data <= "111111";
				when "10100110111001" => data <= "111111";
				when "10100110111010" => data <= "111111";
				when "10100110111011" => data <= "111111";
				when "10100110111100" => data <= "000000";
				when "10100110111101" => data <= "000000";
				when "10100110111110" => data <= "000000";
				when "10100110111111" => data <= "000000";
				when "10100111000000" => data <= "000000";
				when "10100111000001" => data <= "000000";
				when "10100111000010" => data <= "000000";
				when "10100111000011" => data <= "000000";
				when "10100111000100" => data <= "000000";
				when "10100111000101" => data <= "000000";
				when "10100111000110" => data <= "111111";
				when "10100111000111" => data <= "111111";
				when "10100111001000" => data <= "111111";
				when "10100111001001" => data <= "111111";
				when "10100111001010" => data <= "111111";
				when "10100111001011" => data <= "111111";
				when "10100111001100" => data <= "111111";
				when "10100111001101" => data <= "000000";
				when "10100111001110" => data <= "000000";
				when "10100111001111" => data <= "000000";
				when "10100111010000" => data <= "000000";
				when "10100111010001" => data <= "111111";
				when "10100111010010" => data <= "111111";
				when "10100111010011" => data <= "000000";
				when "10100111010100" => data <= "000000";
				when "10100111010101" => data <= "000000";
				when "10100111010110" => data <= "111111";
				when "10100111010111" => data <= "111111";
				when "10100111011000" => data <= "111111";
				when "10100111011001" => data <= "111111";
				when "10100111011010" => data <= "111111";
				when "10100111011011" => data <= "111111";
				when "10100111011100" => data <= "111111";
				when "10100111011101" => data <= "111111";
				when "10100111011110" => data <= "111111";
				when "10100111011111" => data <= "111111";
				when "10100111100000" => data <= "000000";
				when "10100111100001" => data <= "000000";
				when "10100111100010" => data <= "000000";
				when "10100111100011" => data <= "111111";
				when "10100111100100" => data <= "111111";
				when "10100111100101" => data <= "111111";
				when "10100111100110" => data <= "111111";
				when "10100111100111" => data <= "111111";
				when "10100111101000" => data <= "111111";
				when "10100111101001" => data <= "111111";
				when "10100111101010" => data <= "111111";
				when "10100111101011" => data <= "000000";
				when "10100111101100" => data <= "000000";
				when "10100111101101" => data <= "000000";
				when "10100111101110" => data <= "000000";
				when "10100111101111" => data <= "000000";
				when "10100111110000" => data <= "111111";
				when "10100111110001" => data <= "111111";
				when "10100111110010" => data <= "000000";
				when "10100111110011" => data <= "000000";
				when "10100111110100" => data <= "000000";
				when "10100111110101" => data <= "000000";
				when "10100111110110" => data <= "000000";
				when "10100111110111" => data <= "000000";
				when "10100111111000" => data <= "000000";
				when "10100111111001" => data <= "000000";
				when "10100111111010" => data <= "000000";
				when "10100111111011" => data <= "000000";
				when "10100111111100" => data <= "000000";
				when "10100111111101" => data <= "000000";
				when "10100111111110" => data <= "000000";
				when "10100111111111" => data <= "000000";
				when "10101000000000" => data <= "000000";
				when "10101000000001" => data <= "000000";
				when "10101000000010" => data <= "000000";
				when "10101000000011" => data <= "000000";
				when "10101000000100" => data <= "000000";
				when "10101000000101" => data <= "000000";
				when "10101000000110" => data <= "000000";
				when "10101000000111" => data <= "000000";
				when "10101000001000" => data <= "000000";
				when "10101000001001" => data <= "000000";
				when "10101000001010" => data <= "000000";
				when "10101000001011" => data <= "000000";
				when "10101000001100" => data <= "000000";
				when "10101000001101" => data <= "111111";
				when "10101000001110" => data <= "111111";
				when "10101000001111" => data <= "000000";
				when "10101000010000" => data <= "000000";
				when "10101000010001" => data <= "000000";
				when "10101000010010" => data <= "000000";
				when "10101000010011" => data <= "000000";
				when "10101000010100" => data <= "000000";
				when "10101000010101" => data <= "000000";
				when "10101000010110" => data <= "111111";
				when "10101000010111" => data <= "111111";
				when "10101000011000" => data <= "000000";
				when "10101000011001" => data <= "000000";
				when "10101000011010" => data <= "000000";
				when "10101000011011" => data <= "000000";
				when "10101000011100" => data <= "111111";
				when "10101000011101" => data <= "111111";
				when "10101000011110" => data <= "000000";
				when "10101000011111" => data <= "000000";
				when "10101000100000" => data <= "111111";
				when "10101000100001" => data <= "111111";
				when "10101000100010" => data <= "000000";
				when "10101000100011" => data <= "000000";
				when "10101000100100" => data <= "000000";
				when "10101000100101" => data <= "000000";
				when "10101000100110" => data <= "000000";
				when "10101000100111" => data <= "000000";
				when "10101000101000" => data <= "000000";
				when "10101000101001" => data <= "000000";
				when "10101000101010" => data <= "000000";
				when "10101000101011" => data <= "000000";
				when "10101000101100" => data <= "000000";
				when "10101000101101" => data <= "000000";
				when "10101000101110" => data <= "000000";
				when "10101000101111" => data <= "111111";
				when "10101000110000" => data <= "111111";
				when "10101000110001" => data <= "000000";
				when "10101000110010" => data <= "000000";
				when "10101000110011" => data <= "000000";
				when "10101000110100" => data <= "000000";
				when "10101000110101" => data <= "000000";
				when "10101000110110" => data <= "000000";
				when "10101000110111" => data <= "000000";
				when "10101000111000" => data <= "000000";
				when "10101000111001" => data <= "000000";
				when "10101000111010" => data <= "111111";
				when "10101000111011" => data <= "111111";
				when "10101000111100" => data <= "000000";
				when "10101000111101" => data <= "000000";
				when "10101000111110" => data <= "000000";
				when "10101000111111" => data <= "000000";
				when "10101001000000" => data <= "000000";
				when "10101001000001" => data <= "000000";
				when "10101001000010" => data <= "000000";
				when "10101001000011" => data <= "000000";
				when "10101001000100" => data <= "000000";
				when "10101001000101" => data <= "000000";
				when "10101001000110" => data <= "000000";
				when "10101001000111" => data <= "000000";
				when "10101001001000" => data <= "000000";
				when "10101001001001" => data <= "000000";
				when "10101001001010" => data <= "000000";
				when "10101001001011" => data <= "111111";
				when "10101001001100" => data <= "111111";
				when "10101001001101" => data <= "000000";
				when "10101001001110" => data <= "000000";
				when "10101001001111" => data <= "000000";
				when "10101001010000" => data <= "000000";
				when "10101001010001" => data <= "111111";
				when "10101001010010" => data <= "111111";
				when "10101001010011" => data <= "000000";
				when "10101001010100" => data <= "000000";
				when "10101001010101" => data <= "000000";
				when "10101001010110" => data <= "111111";
				when "10101001010111" => data <= "111111";
				when "10101001011000" => data <= "000000";
				when "10101001011001" => data <= "000000";
				when "10101001011010" => data <= "000000";
				when "10101001011011" => data <= "000000";
				when "10101001011100" => data <= "000000";
				when "10101001011101" => data <= "000000";
				when "10101001011110" => data <= "111111";
				when "10101001011111" => data <= "111111";
				when "10101001100000" => data <= "000000";
				when "10101001100001" => data <= "000000";
				when "10101001100010" => data <= "000000";
				when "10101001100011" => data <= "111111";
				when "10101001100100" => data <= "111111";
				when "10101001100101" => data <= "000000";
				when "10101001100110" => data <= "000000";
				when "10101001100111" => data <= "000000";
				when "10101001101000" => data <= "000000";
				when "10101001101001" => data <= "111111";
				when "10101001101010" => data <= "111111";
				when "10101001101011" => data <= "000000";
				when "10101001101100" => data <= "000000";
				when "10101001101101" => data <= "000000";
				when "10101001101110" => data <= "000000";
				when "10101001101111" => data <= "000000";
				when "10101001110000" => data <= "111111";
				when "10101001110001" => data <= "111111";
				when "10101001110010" => data <= "000000";
				when "10101001110011" => data <= "000000";
				when "10101001110100" => data <= "000000";
				when "10101001110101" => data <= "000000";
				when "10101001110110" => data <= "000000";
				when "10101001110111" => data <= "000000";
				when "10101001111000" => data <= "000000";
				when "10101001111001" => data <= "000000";
				when "10101001111010" => data <= "000000";
				when "10101001111011" => data <= "000000";
				when "10101001111100" => data <= "000000";
				when "10101001111101" => data <= "000000";
				when "10101001111110" => data <= "000000";
				when "10101001111111" => data <= "000000";
				when "10101010000000" => data <= "000000";
				when "10101010000001" => data <= "000000";
				when "10101010000010" => data <= "000000";
				when "10101010000011" => data <= "000000";
				when "10101010000100" => data <= "000000";
				when "10101010000101" => data <= "000000";
				when "10101010000110" => data <= "000000";
				when "10101010000111" => data <= "000000";
				when "10101010001000" => data <= "000000";
				when "10101010001001" => data <= "000000";
				when "10101010001010" => data <= "000000";
				when "10101010001011" => data <= "000000";
				when "10101010001100" => data <= "000000";
				when "10101010001101" => data <= "111111";
				when "10101010001110" => data <= "111111";
				when "10101010001111" => data <= "000000";
				when "10101010010000" => data <= "000000";
				when "10101010010001" => data <= "000000";
				when "10101010010010" => data <= "000000";
				when "10101010010011" => data <= "000000";
				when "10101010010100" => data <= "000000";
				when "10101010010101" => data <= "000000";
				when "10101010010110" => data <= "111111";
				when "10101010010111" => data <= "111111";
				when "10101010011000" => data <= "000000";
				when "10101010011001" => data <= "000000";
				when "10101010011010" => data <= "000000";
				when "10101010011011" => data <= "000000";
				when "10101010011100" => data <= "111111";
				when "10101010011101" => data <= "111111";
				when "10101010011110" => data <= "000000";
				when "10101010011111" => data <= "000000";
				when "10101010100000" => data <= "111111";
				when "10101010100001" => data <= "111111";
				when "10101010100010" => data <= "000000";
				when "10101010100011" => data <= "000000";
				when "10101010100100" => data <= "000000";
				when "10101010100101" => data <= "000000";
				when "10101010100110" => data <= "000000";
				when "10101010100111" => data <= "000000";
				when "10101010101000" => data <= "000000";
				when "10101010101001" => data <= "000000";
				when "10101010101010" => data <= "000000";
				when "10101010101011" => data <= "000000";
				when "10101010101100" => data <= "000000";
				when "10101010101101" => data <= "000000";
				when "10101010101110" => data <= "000000";
				when "10101010101111" => data <= "111111";
				when "10101010110000" => data <= "111111";
				when "10101010110001" => data <= "000000";
				when "10101010110010" => data <= "000000";
				when "10101010110011" => data <= "000000";
				when "10101010110100" => data <= "000000";
				when "10101010110101" => data <= "000000";
				when "10101010110110" => data <= "000000";
				when "10101010110111" => data <= "000000";
				when "10101010111000" => data <= "000000";
				when "10101010111001" => data <= "000000";
				when "10101010111010" => data <= "111111";
				when "10101010111011" => data <= "111111";
				when "10101010111100" => data <= "000000";
				when "10101010111101" => data <= "000000";
				when "10101010111110" => data <= "000000";
				when "10101010111111" => data <= "000000";
				when "10101011000000" => data <= "000000";
				when "10101011000001" => data <= "000000";
				when "10101011000010" => data <= "000000";
				when "10101011000011" => data <= "000000";
				when "10101011000100" => data <= "000000";
				when "10101011000101" => data <= "000000";
				when "10101011000110" => data <= "000000";
				when "10101011000111" => data <= "000000";
				when "10101011001000" => data <= "000000";
				when "10101011001001" => data <= "000000";
				when "10101011001010" => data <= "000000";
				when "10101011001011" => data <= "111111";
				when "10101011001100" => data <= "111111";
				when "10101011001101" => data <= "000000";
				when "10101011001110" => data <= "000000";
				when "10101011001111" => data <= "000000";
				when "10101011010000" => data <= "000000";
				when "10101011010001" => data <= "111111";
				when "10101011010010" => data <= "111111";
				when "10101011010011" => data <= "000000";
				when "10101011010100" => data <= "000000";
				when "10101011010101" => data <= "000000";
				when "10101011010110" => data <= "111111";
				when "10101011010111" => data <= "111111";
				when "10101011011000" => data <= "000000";
				when "10101011011001" => data <= "000000";
				when "10101011011010" => data <= "000000";
				when "10101011011011" => data <= "000000";
				when "10101011011100" => data <= "000000";
				when "10101011011101" => data <= "000000";
				when "10101011011110" => data <= "111111";
				when "10101011011111" => data <= "111111";
				when "10101011100000" => data <= "000000";
				when "10101011100001" => data <= "000000";
				when "10101011100010" => data <= "000000";
				when "10101011100011" => data <= "111111";
				when "10101011100100" => data <= "111111";
				when "10101011100101" => data <= "000000";
				when "10101011100110" => data <= "000000";
				when "10101011100111" => data <= "000000";
				when "10101011101000" => data <= "000000";
				when "10101011101001" => data <= "111111";
				when "10101011101010" => data <= "111111";
				when "10101011101011" => data <= "000000";
				when "10101011101100" => data <= "000000";
				when "10101011101101" => data <= "000000";
				when "10101011101110" => data <= "000000";
				when "10101011101111" => data <= "000000";
				when "10101011110000" => data <= "111111";
				when "10101011110001" => data <= "111111";
				when "10101011110010" => data <= "000000";
				when "10101011110011" => data <= "000000";
				when "10101011110100" => data <= "000000";
				when "10101011110101" => data <= "000000";
				when "10101011110110" => data <= "000000";
				when "10101011110111" => data <= "000000";
				when "10101011111000" => data <= "000000";
				when "10101011111001" => data <= "000000";
				when "10101011111010" => data <= "000000";
				when "10101011111011" => data <= "000000";
				when "10101011111100" => data <= "000000";
				when "10101011111101" => data <= "000000";
				when "10101011111110" => data <= "000000";
				when "10101011111111" => data <= "000000";
				when "10101100000000" => data <= "000000";
				when "10101100000001" => data <= "000000";
				when "10101100000010" => data <= "000000";
				when "10101100000011" => data <= "000000";
				when "10101100000100" => data <= "000000";
				when "10101100000101" => data <= "000000";
				when "10101100000110" => data <= "000000";
				when "10101100000111" => data <= "000000";
				when "10101100001000" => data <= "000000";
				when "10101100001001" => data <= "000000";
				when "10101100001010" => data <= "000000";
				when "10101100001011" => data <= "000000";
				when "10101100001100" => data <= "000000";
				when "10101100001101" => data <= "111111";
				when "10101100001110" => data <= "111111";
				when "10101100001111" => data <= "000000";
				when "10101100010000" => data <= "000000";
				when "10101100010001" => data <= "000000";
				when "10101100010010" => data <= "000000";
				when "10101100010011" => data <= "000000";
				when "10101100010100" => data <= "000000";
				when "10101100010101" => data <= "000000";
				when "10101100010110" => data <= "111111";
				when "10101100010111" => data <= "111111";
				when "10101100011000" => data <= "000000";
				when "10101100011001" => data <= "000000";
				when "10101100011010" => data <= "000000";
				when "10101100011011" => data <= "000000";
				when "10101100011100" => data <= "111111";
				when "10101100011101" => data <= "111111";
				when "10101100011110" => data <= "000000";
				when "10101100011111" => data <= "000000";
				when "10101100100000" => data <= "111111";
				when "10101100100001" => data <= "111111";
				when "10101100100010" => data <= "000000";
				when "10101100100011" => data <= "000000";
				when "10101100100100" => data <= "000000";
				when "10101100100101" => data <= "000000";
				when "10101100100110" => data <= "000000";
				when "10101100100111" => data <= "000000";
				when "10101100101000" => data <= "000000";
				when "10101100101001" => data <= "000000";
				when "10101100101010" => data <= "000000";
				when "10101100101011" => data <= "000000";
				when "10101100101100" => data <= "000000";
				when "10101100101101" => data <= "000000";
				when "10101100101110" => data <= "000000";
				when "10101100101111" => data <= "111111";
				when "10101100110000" => data <= "111111";
				when "10101100110001" => data <= "000000";
				when "10101100110010" => data <= "000000";
				when "10101100110011" => data <= "000000";
				when "10101100110100" => data <= "000000";
				when "10101100110101" => data <= "000000";
				when "10101100110110" => data <= "000000";
				when "10101100110111" => data <= "000000";
				when "10101100111000" => data <= "000000";
				when "10101100111001" => data <= "000000";
				when "10101100111010" => data <= "111111";
				when "10101100111011" => data <= "111111";
				when "10101100111100" => data <= "000000";
				when "10101100111101" => data <= "000000";
				when "10101100111110" => data <= "000000";
				when "10101100111111" => data <= "000000";
				when "10101101000000" => data <= "000000";
				when "10101101000001" => data <= "000000";
				when "10101101000010" => data <= "000000";
				when "10101101000011" => data <= "000000";
				when "10101101000100" => data <= "000000";
				when "10101101000101" => data <= "000000";
				when "10101101000110" => data <= "000000";
				when "10101101000111" => data <= "000000";
				when "10101101001000" => data <= "000000";
				when "10101101001001" => data <= "000000";
				when "10101101001010" => data <= "000000";
				when "10101101001011" => data <= "111111";
				when "10101101001100" => data <= "111111";
				when "10101101001101" => data <= "000000";
				when "10101101001110" => data <= "000000";
				when "10101101001111" => data <= "000000";
				when "10101101010000" => data <= "000000";
				when "10101101010001" => data <= "111111";
				when "10101101010010" => data <= "111111";
				when "10101101010011" => data <= "000000";
				when "10101101010100" => data <= "000000";
				when "10101101010101" => data <= "000000";
				when "10101101010110" => data <= "111111";
				when "10101101010111" => data <= "111111";
				when "10101101011000" => data <= "000000";
				when "10101101011001" => data <= "000000";
				when "10101101011010" => data <= "000000";
				when "10101101011011" => data <= "000000";
				when "10101101011100" => data <= "000000";
				when "10101101011101" => data <= "000000";
				when "10101101011110" => data <= "111111";
				when "10101101011111" => data <= "111111";
				when "10101101100000" => data <= "000000";
				when "10101101100001" => data <= "000000";
				when "10101101100010" => data <= "000000";
				when "10101101100011" => data <= "111111";
				when "10101101100100" => data <= "111111";
				when "10101101100101" => data <= "000000";
				when "10101101100110" => data <= "000000";
				when "10101101100111" => data <= "000000";
				when "10101101101000" => data <= "000000";
				when "10101101101001" => data <= "111111";
				when "10101101101010" => data <= "111111";
				when "10101101101011" => data <= "000000";
				when "10101101101100" => data <= "000000";
				when "10101101101101" => data <= "000000";
				when "10101101101110" => data <= "000000";
				when "10101101101111" => data <= "000000";
				when "10101101110000" => data <= "111111";
				when "10101101110001" => data <= "111111";
				when "10101101110010" => data <= "000000";
				when "10101101110011" => data <= "000000";
				when "10101101110100" => data <= "000000";
				when "10101101110101" => data <= "000000";
				when "10101101110110" => data <= "000000";
				when "10101101110111" => data <= "000000";
				when "10101101111000" => data <= "000000";
				when "10101101111001" => data <= "000000";
				when "10101101111010" => data <= "000000";
				when "10101101111011" => data <= "000000";
				when "10101101111100" => data <= "000000";
				when "10101101111101" => data <= "000000";
				when "10101101111110" => data <= "000000";
				when "10101101111111" => data <= "000000";
				when "10101110000000" => data <= "000000";
				when "10101110000001" => data <= "000000";
				when "10101110000010" => data <= "000000";
				when "10101110000011" => data <= "000000";
				when "10101110000100" => data <= "000000";
				when "10101110000101" => data <= "000000";
				when "10101110000110" => data <= "000000";
				when "10101110000111" => data <= "000000";
				when "10101110001000" => data <= "000000";
				when "10101110001001" => data <= "000000";
				when "10101110001010" => data <= "000000";
				when "10101110001011" => data <= "000000";
				when "10101110001100" => data <= "000000";
				when "10101110001101" => data <= "111111";
				when "10101110001110" => data <= "111111";
				when "10101110001111" => data <= "000000";
				when "10101110010000" => data <= "000000";
				when "10101110010001" => data <= "000000";
				when "10101110010010" => data <= "000000";
				when "10101110010011" => data <= "000000";
				when "10101110010100" => data <= "000000";
				when "10101110010101" => data <= "000000";
				when "10101110010110" => data <= "111111";
				when "10101110010111" => data <= "111111";
				when "10101110011000" => data <= "000000";
				when "10101110011001" => data <= "000000";
				when "10101110011010" => data <= "000000";
				when "10101110011011" => data <= "000000";
				when "10101110011100" => data <= "111111";
				when "10101110011101" => data <= "111111";
				when "10101110011110" => data <= "000000";
				when "10101110011111" => data <= "000000";
				when "10101110100000" => data <= "111111";
				when "10101110100001" => data <= "111111";
				when "10101110100010" => data <= "111111";
				when "10101110100011" => data <= "111111";
				when "10101110100100" => data <= "111111";
				when "10101110100101" => data <= "111111";
				when "10101110100110" => data <= "111111";
				when "10101110100111" => data <= "000000";
				when "10101110101000" => data <= "000000";
				when "10101110101001" => data <= "111111";
				when "10101110101010" => data <= "111111";
				when "10101110101011" => data <= "111111";
				when "10101110101100" => data <= "111111";
				when "10101110101101" => data <= "111111";
				when "10101110101110" => data <= "111111";
				when "10101110101111" => data <= "111111";
				when "10101110110000" => data <= "111111";
				when "10101110110001" => data <= "000000";
				when "10101110110010" => data <= "000000";
				when "10101110110011" => data <= "111111";
				when "10101110110100" => data <= "111111";
				when "10101110110101" => data <= "111111";
				when "10101110110110" => data <= "111111";
				when "10101110110111" => data <= "111111";
				when "10101110111000" => data <= "111111";
				when "10101110111001" => data <= "111111";
				when "10101110111010" => data <= "111111";
				when "10101110111011" => data <= "111111";
				when "10101110111100" => data <= "000000";
				when "10101110111101" => data <= "000000";
				when "10101110111110" => data <= "000000";
				when "10101110111111" => data <= "000000";
				when "10101111000000" => data <= "000000";
				when "10101111000001" => data <= "000000";
				when "10101111000010" => data <= "000000";
				when "10101111000011" => data <= "000000";
				when "10101111000100" => data <= "111111";
				when "10101111000101" => data <= "111111";
				when "10101111000110" => data <= "111111";
				when "10101111000111" => data <= "111111";
				when "10101111001000" => data <= "111111";
				when "10101111001001" => data <= "111111";
				when "10101111001010" => data <= "111111";
				when "10101111001011" => data <= "111111";
				when "10101111001100" => data <= "111111";
				when "10101111001101" => data <= "000000";
				when "10101111001110" => data <= "000000";
				when "10101111001111" => data <= "000000";
				when "10101111010000" => data <= "000000";
				when "10101111010001" => data <= "111111";
				when "10101111010010" => data <= "111111";
				when "10101111010011" => data <= "000000";
				when "10101111010100" => data <= "000000";
				when "10101111010101" => data <= "000000";
				when "10101111010110" => data <= "111111";
				when "10101111010111" => data <= "111111";
				when "10101111011000" => data <= "000000";
				when "10101111011001" => data <= "000000";
				when "10101111011010" => data <= "000000";
				when "10101111011011" => data <= "000000";
				when "10101111011100" => data <= "000000";
				when "10101111011101" => data <= "000000";
				when "10101111011110" => data <= "111111";
				when "10101111011111" => data <= "111111";
				when "10101111100000" => data <= "000000";
				when "10101111100001" => data <= "000000";
				when "10101111100010" => data <= "000000";
				when "10101111100011" => data <= "111111";
				when "10101111100100" => data <= "111111";
				when "10101111100101" => data <= "000000";
				when "10101111100110" => data <= "000000";
				when "10101111100111" => data <= "000000";
				when "10101111101000" => data <= "000000";
				when "10101111101001" => data <= "111111";
				when "10101111101010" => data <= "111111";
				when "10101111101011" => data <= "000000";
				when "10101111101100" => data <= "000000";
				when "10101111101101" => data <= "000000";
				when "10101111101110" => data <= "000000";
				when "10101111101111" => data <= "000000";
				when "10101111110000" => data <= "111111";
				when "10101111110001" => data <= "111111";
				when "10101111110010" => data <= "000000";
				when "10101111110011" => data <= "000000";
				when "10101111110100" => data <= "000000";
				when "10101111110101" => data <= "000000";
				when "10101111110110" => data <= "000000";
				when "10101111110111" => data <= "000000";
				when "10101111111000" => data <= "000000";
				when "10101111111001" => data <= "000000";
				when "10101111111010" => data <= "000000";
				when "10101111111011" => data <= "000000";
				when "10101111111100" => data <= "000000";
				when "10101111111101" => data <= "000000";
				when "10101111111110" => data <= "000000";
				when "10101111111111" => data <= "000000";
				when "10110000000000" => data <= "000000";
				when "10110000000001" => data <= "000000";
				when "10110000000010" => data <= "000000";
				when "10110000000011" => data <= "000000";
				when "10110000000100" => data <= "000000";
				when "10110000000101" => data <= "000000";
				when "10110000000110" => data <= "000000";
				when "10110000000111" => data <= "000000";
				when "10110000001000" => data <= "000000";
				when "10110000001001" => data <= "000000";
				when "10110000001010" => data <= "000000";
				when "10110000001011" => data <= "000000";
				when "10110000001100" => data <= "000000";
				when "10110000001101" => data <= "111111";
				when "10110000001110" => data <= "111111";
				when "10110000001111" => data <= "000000";
				when "10110000010000" => data <= "000000";
				when "10110000010001" => data <= "000000";
				when "10110000010010" => data <= "000000";
				when "10110000010011" => data <= "000000";
				when "10110000010100" => data <= "000000";
				when "10110000010101" => data <= "000000";
				when "10110000010110" => data <= "111111";
				when "10110000010111" => data <= "111111";
				when "10110000011000" => data <= "000000";
				when "10110000011001" => data <= "000000";
				when "10110000011010" => data <= "000000";
				when "10110000011011" => data <= "000000";
				when "10110000011100" => data <= "111111";
				when "10110000011101" => data <= "111111";
				when "10110000011110" => data <= "000000";
				when "10110000011111" => data <= "000000";
				when "10110000100000" => data <= "111111";
				when "10110000100001" => data <= "111111";
				when "10110000100010" => data <= "111111";
				when "10110000100011" => data <= "111111";
				when "10110000100100" => data <= "111111";
				when "10110000100101" => data <= "111111";
				when "10110000100110" => data <= "111111";
				when "10110000100111" => data <= "000000";
				when "10110000101000" => data <= "000000";
				when "10110000101001" => data <= "111111";
				when "10110000101010" => data <= "111111";
				when "10110000101011" => data <= "111111";
				when "10110000101100" => data <= "111111";
				when "10110000101101" => data <= "111111";
				when "10110000101110" => data <= "111111";
				when "10110000101111" => data <= "000000";
				when "10110000110000" => data <= "000000";
				when "10110000110001" => data <= "000000";
				when "10110000110010" => data <= "000000";
				when "10110000110011" => data <= "111111";
				when "10110000110100" => data <= "111111";
				when "10110000110101" => data <= "111111";
				when "10110000110110" => data <= "111111";
				when "10110000110111" => data <= "111111";
				when "10110000111000" => data <= "111111";
				when "10110000111001" => data <= "111111";
				when "10110000111010" => data <= "000000";
				when "10110000111011" => data <= "000000";
				when "10110000111100" => data <= "000000";
				when "10110000111101" => data <= "000000";
				when "10110000111110" => data <= "000000";
				when "10110000111111" => data <= "000000";
				when "10110001000000" => data <= "000000";
				when "10110001000001" => data <= "000000";
				when "10110001000010" => data <= "000000";
				when "10110001000011" => data <= "000000";
				when "10110001000100" => data <= "111111";
				when "10110001000101" => data <= "111111";
				when "10110001000110" => data <= "111111";
				when "10110001000111" => data <= "111111";
				when "10110001001000" => data <= "111111";
				when "10110001001001" => data <= "111111";
				when "10110001001010" => data <= "111111";
				when "10110001001011" => data <= "000000";
				when "10110001001100" => data <= "000000";
				when "10110001001101" => data <= "000000";
				when "10110001001110" => data <= "000000";
				when "10110001001111" => data <= "000000";
				when "10110001010000" => data <= "000000";
				when "10110001010001" => data <= "111111";
				when "10110001010010" => data <= "111111";
				when "10110001010011" => data <= "000000";
				when "10110001010100" => data <= "000000";
				when "10110001010101" => data <= "000000";
				when "10110001010110" => data <= "111111";
				when "10110001010111" => data <= "111111";
				when "10110001011000" => data <= "000000";
				when "10110001011001" => data <= "000000";
				when "10110001011010" => data <= "000000";
				when "10110001011011" => data <= "000000";
				when "10110001011100" => data <= "000000";
				when "10110001011101" => data <= "000000";
				when "10110001011110" => data <= "111111";
				when "10110001011111" => data <= "111111";
				when "10110001100000" => data <= "000000";
				when "10110001100001" => data <= "000000";
				when "10110001100010" => data <= "000000";
				when "10110001100011" => data <= "111111";
				when "10110001100100" => data <= "111111";
				when "10110001100101" => data <= "000000";
				when "10110001100110" => data <= "000000";
				when "10110001100111" => data <= "000000";
				when "10110001101000" => data <= "000000";
				when "10110001101001" => data <= "111111";
				when "10110001101010" => data <= "111111";
				when "10110001101011" => data <= "000000";
				when "10110001101100" => data <= "000000";
				when "10110001101101" => data <= "000000";
				when "10110001101110" => data <= "000000";
				when "10110001101111" => data <= "000000";
				when "10110001110000" => data <= "111111";
				when "10110001110001" => data <= "111111";
				when "10110001110010" => data <= "000000";
				when "10110001110011" => data <= "000000";
				when "10110001110100" => data <= "000000";
				when "10110001110101" => data <= "000000";
				when "10110001110110" => data <= "000000";
				when "10110001110111" => data <= "000000";
				when "10110001111000" => data <= "000000";
				when "10110001111001" => data <= "000000";
				when "10110001111010" => data <= "000000";
				when "10110001111011" => data <= "000000";
				when "10110001111100" => data <= "000000";
				when "10110001111101" => data <= "000000";
				when "10110001111110" => data <= "000000";
				when "10110001111111" => data <= "000000";
				when "10110010000000" => data <= "000000";
				when "10110010000001" => data <= "000000";
				when "10110010000010" => data <= "000000";
				when "10110010000011" => data <= "000000";
				when "10110010000100" => data <= "000000";
				when "10110010000101" => data <= "000000";
				when "10110010000110" => data <= "000000";
				when "10110010000111" => data <= "000000";
				when "10110010001000" => data <= "000000";
				when "10110010001001" => data <= "000000";
				when "10110010001010" => data <= "000000";
				when "10110010001011" => data <= "000000";
				when "10110010001100" => data <= "000000";
				when "10110010001101" => data <= "000000";
				when "10110010001110" => data <= "000000";
				when "10110010001111" => data <= "000000";
				when "10110010010000" => data <= "000000";
				when "10110010010001" => data <= "000000";
				when "10110010010010" => data <= "000000";
				when "10110010010011" => data <= "000000";
				when "10110010010100" => data <= "000000";
				when "10110010010101" => data <= "000000";
				when "10110010010110" => data <= "000000";
				when "10110010010111" => data <= "000000";
				when "10110010011000" => data <= "000000";
				when "10110010011001" => data <= "000000";
				when "10110010011010" => data <= "000000";
				when "10110010011011" => data <= "000000";
				when "10110010011100" => data <= "000000";
				when "10110010011101" => data <= "000000";
				when "10110010011110" => data <= "000000";
				when "10110010011111" => data <= "000000";
				when "10110010100000" => data <= "000000";
				when "10110010100001" => data <= "000000";
				when "10110010100010" => data <= "000000";
				when "10110010100011" => data <= "000000";
				when "10110010100100" => data <= "000000";
				when "10110010100101" => data <= "000000";
				when "10110010100110" => data <= "000000";
				when "10110010100111" => data <= "000000";
				when "10110010101000" => data <= "000000";
				when "10110010101001" => data <= "000000";
				when "10110010101010" => data <= "000000";
				when "10110010101011" => data <= "000000";
				when "10110010101100" => data <= "000000";
				when "10110010101101" => data <= "000000";
				when "10110010101110" => data <= "000000";
				when "10110010101111" => data <= "000000";
				when "10110010110000" => data <= "000000";
				when "10110010110001" => data <= "000000";
				when "10110010110010" => data <= "000000";
				when "10110010110011" => data <= "000000";
				when "10110010110100" => data <= "000000";
				when "10110010110101" => data <= "000000";
				when "10110010110110" => data <= "000000";
				when "10110010110111" => data <= "000000";
				when "10110010111000" => data <= "000000";
				when "10110010111001" => data <= "000000";
				when "10110010111010" => data <= "000000";
				when "10110010111011" => data <= "000000";
				when "10110010111100" => data <= "000000";
				when "10110010111101" => data <= "000000";
				when "10110010111110" => data <= "000000";
				when "10110010111111" => data <= "000000";
				when "10110011000000" => data <= "000000";
				when "10110011000001" => data <= "000000";
				when "10110011000010" => data <= "000000";
				when "10110011000011" => data <= "000000";
				when "10110011000100" => data <= "000000";
				when "10110011000101" => data <= "000000";
				when "10110011000110" => data <= "000000";
				when "10110011000111" => data <= "000000";
				when "10110011001000" => data <= "000000";
				when "10110011001001" => data <= "000000";
				when "10110011001010" => data <= "000000";
				when "10110011001011" => data <= "000000";
				when "10110011001100" => data <= "000000";
				when "10110011001101" => data <= "000000";
				when "10110011001110" => data <= "000000";
				when "10110011001111" => data <= "000000";
				when "10110011010000" => data <= "000000";
				when "10110011010001" => data <= "000000";
				when "10110011010010" => data <= "000000";
				when "10110011010011" => data <= "000000";
				when "10110011010100" => data <= "000000";
				when "10110011010101" => data <= "000000";
				when "10110011010110" => data <= "000000";
				when "10110011010111" => data <= "000000";
				when "10110011011000" => data <= "000000";
				when "10110011011001" => data <= "000000";
				when "10110011011010" => data <= "000000";
				when "10110011011011" => data <= "000000";
				when "10110011011100" => data <= "000000";
				when "10110011011101" => data <= "000000";
				when "10110011011110" => data <= "000000";
				when "10110011011111" => data <= "000000";
				when "10110011100000" => data <= "000000";
				when "10110011100001" => data <= "000000";
				when "10110011100010" => data <= "000000";
				when "10110011100011" => data <= "000000";
				when "10110011100100" => data <= "000000";
				when "10110011100101" => data <= "000000";
				when "10110011100110" => data <= "000000";
				when "10110011100111" => data <= "000000";
				when "10110011101000" => data <= "000000";
				when "10110011101001" => data <= "000000";
				when "10110011101010" => data <= "000000";
				when "10110011101011" => data <= "000000";
				when "10110011101100" => data <= "000000";
				when "10110011101101" => data <= "000000";
				when "10110011101110" => data <= "000000";
				when "10110011101111" => data <= "000000";
				when "10110011110000" => data <= "000000";
				when "10110011110001" => data <= "000000";
				when "10110011110010" => data <= "000000";
				when "10110011110011" => data <= "000000";
				when "10110011110100" => data <= "000000";
				when "10110011110101" => data <= "000000";
				when "10110011110110" => data <= "000000";
				when "10110011110111" => data <= "000000";
				when "10110011111000" => data <= "000000";
				when "10110011111001" => data <= "000000";
				when "10110011111010" => data <= "000000";
				when "10110011111011" => data <= "000000";
				when "10110011111100" => data <= "000000";
				when "10110011111101" => data <= "000000";
				when "10110011111110" => data <= "000000";
				when "10110011111111" => data <= "000000";
				when "10110100000000" => data <= "000000";
				when "10110100000001" => data <= "000000";
				when "10110100000010" => data <= "000000";
				when "10110100000011" => data <= "000000";
				when "10110100000100" => data <= "000000";
				when "10110100000101" => data <= "000000";
				when "10110100000110" => data <= "000000";
				when "10110100000111" => data <= "000000";
				when "10110100001000" => data <= "000000";
				when "10110100001001" => data <= "000000";
				when "10110100001010" => data <= "000000";
				when "10110100001011" => data <= "000000";
				when "10110100001100" => data <= "000000";
				when "10110100001101" => data <= "000000";
				when "10110100001110" => data <= "000000";
				when "10110100001111" => data <= "000000";
				when "10110100010000" => data <= "000000";
				when "10110100010001" => data <= "000000";
				when "10110100010010" => data <= "000000";
				when "10110100010011" => data <= "000000";
				when "10110100010100" => data <= "000000";
				when "10110100010101" => data <= "000000";
				when "10110100010110" => data <= "000000";
				when "10110100010111" => data <= "000000";
				when "10110100011000" => data <= "000000";
				when "10110100011001" => data <= "000000";
				when "10110100011010" => data <= "000000";
				when "10110100011011" => data <= "000000";
				when "10110100011100" => data <= "000000";
				when "10110100011101" => data <= "000000";
				when "10110100011110" => data <= "000000";
				when "10110100011111" => data <= "000000";
				when "10110100100000" => data <= "000000";
				when "10110100100001" => data <= "000000";
				when "10110100100010" => data <= "000000";
				when "10110100100011" => data <= "000000";
				when "10110100100100" => data <= "000000";
				when "10110100100101" => data <= "000000";
				when "10110100100110" => data <= "000000";
				when "10110100100111" => data <= "000000";
				when "10110100101000" => data <= "000000";
				when "10110100101001" => data <= "000000";
				when "10110100101010" => data <= "000000";
				when "10110100101011" => data <= "000000";
				when "10110100101100" => data <= "000000";
				when "10110100101101" => data <= "000000";
				when "10110100101110" => data <= "000000";
				when "10110100101111" => data <= "000000";
				when "10110100110000" => data <= "000000";
				when "10110100110001" => data <= "000000";
				when "10110100110010" => data <= "000000";
				when "10110100110011" => data <= "000000";
				when "10110100110100" => data <= "000000";
				when "10110100110101" => data <= "000000";
				when "10110100110110" => data <= "000000";
				when "10110100110111" => data <= "000000";
				when "10110100111000" => data <= "000000";
				when "10110100111001" => data <= "000000";
				when "10110100111010" => data <= "000000";
				when "10110100111011" => data <= "000000";
				when "10110100111100" => data <= "000000";
				when "10110100111101" => data <= "000000";
				when "10110100111110" => data <= "000000";
				when "10110100111111" => data <= "000000";
				when "10110101000000" => data <= "000000";
				when "10110101000001" => data <= "000000";
				when "10110101000010" => data <= "000000";
				when "10110101000011" => data <= "000000";
				when "10110101000100" => data <= "000000";
				when "10110101000101" => data <= "000000";
				when "10110101000110" => data <= "000000";
				when "10110101000111" => data <= "000000";
				when "10110101001000" => data <= "000000";
				when "10110101001001" => data <= "000000";
				when "10110101001010" => data <= "000000";
				when "10110101001011" => data <= "000000";
				when "10110101001100" => data <= "000000";
				when "10110101001101" => data <= "000000";
				when "10110101001110" => data <= "000000";
				when "10110101001111" => data <= "000000";
				when "10110101010000" => data <= "000000";
				when "10110101010001" => data <= "000000";
				when "10110101010010" => data <= "000000";
				when "10110101010011" => data <= "000000";
				when "10110101010100" => data <= "000000";
				when "10110101010101" => data <= "000000";
				when "10110101010110" => data <= "000000";
				when "10110101010111" => data <= "000000";
				when "10110101011000" => data <= "000000";
				when "10110101011001" => data <= "000000";
				when "10110101011010" => data <= "000000";
				when "10110101011011" => data <= "000000";
				when "10110101011100" => data <= "000000";
				when "10110101011101" => data <= "000000";
				when "10110101011110" => data <= "000000";
				when "10110101011111" => data <= "000000";
				when "10110101100000" => data <= "000000";
				when "10110101100001" => data <= "000000";
				when "10110101100010" => data <= "000000";
				when "10110101100011" => data <= "000000";
				when "10110101100100" => data <= "000000";
				when "10110101100101" => data <= "000000";
				when "10110101100110" => data <= "000000";
				when "10110101100111" => data <= "000000";
				when "10110101101000" => data <= "000000";
				when "10110101101001" => data <= "000000";
				when "10110101101010" => data <= "000000";
				when "10110101101011" => data <= "000000";
				when "10110101101100" => data <= "000000";
				when "10110101101101" => data <= "000000";
				when "10110101101110" => data <= "000000";
				when "10110101101111" => data <= "000000";
				when "10110101110000" => data <= "000000";
				when "10110101110001" => data <= "000000";
				when "10110101110010" => data <= "000000";
				when "10110101110011" => data <= "000000";
				when "10110101110100" => data <= "000000";
				when "10110101110101" => data <= "000000";
				when "10110101110110" => data <= "000000";
				when "10110101110111" => data <= "000000";
				when "10110101111000" => data <= "000000";
				when "10110101111001" => data <= "000000";
				when "10110101111010" => data <= "000000";
				when "10110101111011" => data <= "000000";
				when "10110101111100" => data <= "000000";
				when "10110101111101" => data <= "000000";
				when "10110101111110" => data <= "000000";
				when "10110101111111" => data <= "000000";
				when "10110110000000" => data <= "000000";
				when "10110110000001" => data <= "000000";
				when "10110110000010" => data <= "000000";
				when "10110110000011" => data <= "000000";
				when "10110110000100" => data <= "000000";
				when "10110110000101" => data <= "000000";
				when "10110110000110" => data <= "000000";
				when "10110110000111" => data <= "000000";
				when "10110110001000" => data <= "000000";
				when "10110110001001" => data <= "000000";
				when "10110110001010" => data <= "000000";
				when "10110110001011" => data <= "000000";
				when "10110110001100" => data <= "000000";
				when "10110110001101" => data <= "000000";
				when "10110110001110" => data <= "000000";
				when "10110110001111" => data <= "000000";
				when "10110110010000" => data <= "000000";
				when "10110110010001" => data <= "000000";
				when "10110110010010" => data <= "000000";
				when "10110110010011" => data <= "000000";
				when "10110110010100" => data <= "000000";
				when "10110110010101" => data <= "000000";
				when "10110110010110" => data <= "000000";
				when "10110110010111" => data <= "000000";
				when "10110110011000" => data <= "000000";
				when "10110110011001" => data <= "000000";
				when "10110110011010" => data <= "000000";
				when "10110110011011" => data <= "000000";
				when "10110110011100" => data <= "000000";
				when "10110110011101" => data <= "000000";
				when "10110110011110" => data <= "000000";
				when "10110110011111" => data <= "000000";
				when "10110110100000" => data <= "000000";
				when "10110110100001" => data <= "000000";
				when "10110110100010" => data <= "000000";
				when "10110110100011" => data <= "000000";
				when "10110110100100" => data <= "000000";
				when "10110110100101" => data <= "000000";
				when "10110110100110" => data <= "000000";
				when "10110110100111" => data <= "000000";
				when "10110110101000" => data <= "000000";
				when "10110110101001" => data <= "000000";
				when "10110110101010" => data <= "000000";
				when "10110110101011" => data <= "000000";
				when "10110110101100" => data <= "000000";
				when "10110110101101" => data <= "000000";
				when "10110110101110" => data <= "000000";
				when "10110110101111" => data <= "000000";
				when "10110110110000" => data <= "000000";
				when "10110110110001" => data <= "000000";
				when "10110110110010" => data <= "000000";
				when "10110110110011" => data <= "000000";
				when "10110110110100" => data <= "000000";
				when "10110110110101" => data <= "000000";
				when "10110110110110" => data <= "000000";
				when "10110110110111" => data <= "000000";
				when "10110110111000" => data <= "000000";
				when "10110110111001" => data <= "000000";
				when "10110110111010" => data <= "000000";
				when "10110110111011" => data <= "000000";
				when "10110110111100" => data <= "000000";
				when "10110110111101" => data <= "000000";
				when "10110110111110" => data <= "000000";
				when "10110110111111" => data <= "000000";
				when "10110111000000" => data <= "000000";
				when "10110111000001" => data <= "000000";
				when "10110111000010" => data <= "000000";
				when "10110111000011" => data <= "000000";
				when "10110111000100" => data <= "000000";
				when "10110111000101" => data <= "000000";
				when "10110111000110" => data <= "000000";
				when "10110111000111" => data <= "000000";
				when "10110111001000" => data <= "000000";
				when "10110111001001" => data <= "000000";
				when "10110111001010" => data <= "000000";
				when "10110111001011" => data <= "000000";
				when "10110111001100" => data <= "000000";
				when "10110111001101" => data <= "000000";
				when "10110111001110" => data <= "000000";
				when "10110111001111" => data <= "000000";
				when "10110111010000" => data <= "000000";
				when "10110111010001" => data <= "000000";
				when "10110111010010" => data <= "000000";
				when "10110111010011" => data <= "000000";
				when "10110111010100" => data <= "000000";
				when "10110111010101" => data <= "000000";
				when "10110111010110" => data <= "000000";
				when "10110111010111" => data <= "000000";
				when "10110111011000" => data <= "000000";
				when "10110111011001" => data <= "000000";
				when "10110111011010" => data <= "000000";
				when "10110111011011" => data <= "000000";
				when "10110111011100" => data <= "000000";
				when "10110111011101" => data <= "000000";
				when "10110111011110" => data <= "000000";
				when "10110111011111" => data <= "000000";
				when "10110111100000" => data <= "000000";
				when "10110111100001" => data <= "000000";
				when "10110111100010" => data <= "000000";
				when "10110111100011" => data <= "000000";
				when "10110111100100" => data <= "000000";
				when "10110111100101" => data <= "000000";
				when "10110111100110" => data <= "000000";
				when "10110111100111" => data <= "000000";
				when "10110111101000" => data <= "000000";
				when "10110111101001" => data <= "000000";
				when "10110111101010" => data <= "000000";
				when "10110111101011" => data <= "000000";
				when "10110111101100" => data <= "000000";
				when "10110111101101" => data <= "000000";
				when "10110111101110" => data <= "000000";
				when "10110111101111" => data <= "000000";
				when "10110111110000" => data <= "000000";
				when "10110111110001" => data <= "000000";
				when "10110111110010" => data <= "000000";
				when "10110111110011" => data <= "000000";
				when "10110111110100" => data <= "000000";
				when "10110111110101" => data <= "000000";
				when "10110111110110" => data <= "000000";
				when "10110111110111" => data <= "000000";
				when "10110111111000" => data <= "000000";
				when "10110111111001" => data <= "000000";
				when "10110111111010" => data <= "000000";
				when "10110111111011" => data <= "000000";
				when "10110111111100" => data <= "000000";
				when "10110111111101" => data <= "000000";
				when "10110111111110" => data <= "000000";
				when "10110111111111" => data <= "000000";
				when "10111000000000" => data <= "000000";
				when "10111000000001" => data <= "000000";
				when "10111000000010" => data <= "000000";
				when "10111000000011" => data <= "000000";
				when "10111000000100" => data <= "000000";
				when "10111000000101" => data <= "000000";
				when "10111000000110" => data <= "000000";
				when "10111000000111" => data <= "000000";
				when "10111000001000" => data <= "000000";
				when "10111000001001" => data <= "000000";
				when "10111000001010" => data <= "000000";
				when "10111000001011" => data <= "000000";
				when "10111000001100" => data <= "000000";
				when "10111000001101" => data <= "000000";
				when "10111000001110" => data <= "000000";
				when "10111000001111" => data <= "000000";
				when "10111000010000" => data <= "000000";
				when "10111000010001" => data <= "000000";
				when "10111000010010" => data <= "000000";
				when "10111000010011" => data <= "000000";
				when "10111000010100" => data <= "000000";
				when "10111000010101" => data <= "000000";
				when "10111000010110" => data <= "000000";
				when "10111000010111" => data <= "000000";
				when "10111000011000" => data <= "000000";
				when "10111000011001" => data <= "000000";
				when "10111000011010" => data <= "000000";
				when "10111000011011" => data <= "000000";
				when "10111000011100" => data <= "000000";
				when "10111000011101" => data <= "000000";
				when "10111000011110" => data <= "000000";
				when "10111000011111" => data <= "000000";
				when "10111000100000" => data <= "000000";
				when "10111000100001" => data <= "000000";
				when "10111000100010" => data <= "000000";
				when "10111000100011" => data <= "000000";
				when "10111000100100" => data <= "000000";
				when "10111000100101" => data <= "000000";
				when "10111000100110" => data <= "000000";
				when "10111000100111" => data <= "000000";
				when "10111000101000" => data <= "000000";
				when "10111000101001" => data <= "000000";
				when "10111000101010" => data <= "000000";
				when "10111000101011" => data <= "000000";
				when "10111000101100" => data <= "000000";
				when "10111000101101" => data <= "000000";
				when "10111000101110" => data <= "000000";
				when "10111000101111" => data <= "000000";
				when "10111000110000" => data <= "000000";
				when "10111000110001" => data <= "000000";
				when "10111000110010" => data <= "000000";
				when "10111000110011" => data <= "000000";
				when "10111000110100" => data <= "000000";
				when "10111000110101" => data <= "000000";
				when "10111000110110" => data <= "000000";
				when "10111000110111" => data <= "000000";
				when "10111000111000" => data <= "000000";
				when "10111000111001" => data <= "000000";
				when "10111000111010" => data <= "000000";
				when "10111000111011" => data <= "000000";
				when "10111000111100" => data <= "000000";
				when "10111000111101" => data <= "000000";
				when "10111000111110" => data <= "000000";
				when "10111000111111" => data <= "000000";
				when "10111001000000" => data <= "000000";
				when "10111001000001" => data <= "000000";
				when "10111001000010" => data <= "000000";
				when "10111001000011" => data <= "000000";
				when "10111001000100" => data <= "000000";
				when "10111001000101" => data <= "000000";
				when "10111001000110" => data <= "000000";
				when "10111001000111" => data <= "000000";
				when "10111001001000" => data <= "000000";
				when "10111001001001" => data <= "000000";
				when "10111001001010" => data <= "000000";
				when "10111001001011" => data <= "000000";
				when "10111001001100" => data <= "000000";
				when "10111001001101" => data <= "000000";
				when "10111001001110" => data <= "000000";
				when "10111001001111" => data <= "000000";
				when "10111001010000" => data <= "000000";
				when "10111001010001" => data <= "000000";
				when "10111001010010" => data <= "000000";
				when "10111001010011" => data <= "000000";
				when "10111001010100" => data <= "000000";
				when "10111001010101" => data <= "000000";
				when "10111001010110" => data <= "000000";
				when "10111001010111" => data <= "000000";
				when "10111001011000" => data <= "000000";
				when "10111001011001" => data <= "000000";
				when "10111001011010" => data <= "000000";
				when "10111001011011" => data <= "000000";
				when "10111001011100" => data <= "000000";
				when "10111001011101" => data <= "000000";
				when "10111001011110" => data <= "000000";
				when "10111001011111" => data <= "000000";
				when "10111001100000" => data <= "000000";
				when "10111001100001" => data <= "000000";
				when "10111001100010" => data <= "000000";
				when "10111001100011" => data <= "000000";
				when "10111001100100" => data <= "000000";
				when "10111001100101" => data <= "000000";
				when "10111001100110" => data <= "000000";
				when "10111001100111" => data <= "000000";
				when "10111001101000" => data <= "000000";
				when "10111001101001" => data <= "000000";
				when "10111001101010" => data <= "000000";
				when "10111001101011" => data <= "000000";
				when "10111001101100" => data <= "000000";
				when "10111001101101" => data <= "000000";
				when "10111001101110" => data <= "000000";
				when "10111001101111" => data <= "000000";
				when "10111001110000" => data <= "000000";
				when "10111001110001" => data <= "000000";
				when "10111001110010" => data <= "000000";
				when "10111001110011" => data <= "000000";
				when "10111001110100" => data <= "000000";
				when "10111001110101" => data <= "000000";
				when "10111001110110" => data <= "000000";
				when "10111001110111" => data <= "000000";
				when "10111001111000" => data <= "000000";
				when "10111001111001" => data <= "000000";
				when "10111001111010" => data <= "000000";
				when "10111001111011" => data <= "000000";
				when "10111001111100" => data <= "000000";
				when "10111001111101" => data <= "000000";
				when "10111001111110" => data <= "000000";
				when "10111001111111" => data <= "000000";
				when "10111010000000" => data <= "000000";
				when "10111010000001" => data <= "000000";
				when "10111010000010" => data <= "000000";
				when "10111010000011" => data <= "000000";
				when "10111010000100" => data <= "000000";
				when "10111010000101" => data <= "000000";
				when "10111010000110" => data <= "000000";
				when "10111010000111" => data <= "000000";
				when "10111010001000" => data <= "000000";
				when "10111010001001" => data <= "000000";
				when "10111010001010" => data <= "000000";
				when "10111010001011" => data <= "000000";
				when "10111010001100" => data <= "000000";
				when "10111010001101" => data <= "000000";
				when "10111010001110" => data <= "000000";
				when "10111010001111" => data <= "000000";
				when "10111010010000" => data <= "000000";
				when "10111010010001" => data <= "000000";
				when "10111010010010" => data <= "000000";
				when "10111010010011" => data <= "000000";
				when "10111010010100" => data <= "000000";
				when "10111010010101" => data <= "000000";
				when "10111010010110" => data <= "000000";
				when "10111010010111" => data <= "000000";
				when "10111010011000" => data <= "000000";
				when "10111010011001" => data <= "000000";
				when "10111010011010" => data <= "000000";
				when "10111010011011" => data <= "000000";
				when "10111010011100" => data <= "000000";
				when "10111010011101" => data <= "000000";
				when "10111010011110" => data <= "000000";
				when "10111010011111" => data <= "000000";
				when "10111010100000" => data <= "000000";
				when "10111010100001" => data <= "000000";
				when "10111010100010" => data <= "000000";
				when "10111010100011" => data <= "000000";
				when "10111010100100" => data <= "000000";
				when "10111010100101" => data <= "000000";
				when "10111010100110" => data <= "000000";
				when "10111010100111" => data <= "000000";
				when "10111010101000" => data <= "000000";
				when "10111010101001" => data <= "000000";
				when "10111010101010" => data <= "000000";
				when "10111010101011" => data <= "000000";
				when "10111010101100" => data <= "000000";
				when "10111010101101" => data <= "000000";
				when "10111010101110" => data <= "000000";
				when "10111010101111" => data <= "000000";
				when "10111010110000" => data <= "000000";
				when "10111010110001" => data <= "000000";
				when "10111010110010" => data <= "000000";
				when "10111010110011" => data <= "000000";
				when "10111010110100" => data <= "000000";
				when "10111010110101" => data <= "000000";
				when "10111010110110" => data <= "000000";
				when "10111010110111" => data <= "000000";
				when "10111010111000" => data <= "000000";
				when "10111010111001" => data <= "000000";
				when "10111010111010" => data <= "000000";
				when "10111010111011" => data <= "000000";
				when "10111010111100" => data <= "000000";
				when "10111010111101" => data <= "000000";
				when "10111010111110" => data <= "000000";
				when "10111010111111" => data <= "000000";
				when "10111011000000" => data <= "000000";
				when "10111011000001" => data <= "000000";
				when "10111011000010" => data <= "000000";
				when "10111011000011" => data <= "000000";
				when "10111011000100" => data <= "000000";
				when "10111011000101" => data <= "000000";
				when "10111011000110" => data <= "000000";
				when "10111011000111" => data <= "000000";
				when "10111011001000" => data <= "000000";
				when "10111011001001" => data <= "000000";
				when "10111011001010" => data <= "000000";
				when "10111011001011" => data <= "000000";
				when "10111011001100" => data <= "000000";
				when "10111011001101" => data <= "000000";
				when "10111011001110" => data <= "000000";
				when "10111011001111" => data <= "000000";
				when "10111011010000" => data <= "000000";
				when "10111011010001" => data <= "000000";
				when "10111011010010" => data <= "000000";
				when "10111011010011" => data <= "000000";
				when "10111011010100" => data <= "000000";
				when "10111011010101" => data <= "000000";
				when "10111011010110" => data <= "000000";
				when "10111011010111" => data <= "000000";
				when "10111011011000" => data <= "000000";
				when "10111011011001" => data <= "000000";
				when "10111011011010" => data <= "000000";
				when "10111011011011" => data <= "000000";
				when "10111011011100" => data <= "000000";
				when "10111011011101" => data <= "000000";
				when "10111011011110" => data <= "000000";
				when "10111011011111" => data <= "000000";
				when "10111011100000" => data <= "000000";
				when "10111011100001" => data <= "000000";
				when "10111011100010" => data <= "000000";
				when "10111011100011" => data <= "000000";
				when "10111011100100" => data <= "000000";
				when "10111011100101" => data <= "000000";
				when "10111011100110" => data <= "000000";
				when "10111011100111" => data <= "000000";
				when "10111011101000" => data <= "000000";
				when "10111011101001" => data <= "000000";
				when "10111011101010" => data <= "000000";
				when "10111011101011" => data <= "000000";
				when "10111011101100" => data <= "000000";
				when "10111011101101" => data <= "000000";
				when "10111011101110" => data <= "000000";
				when "10111011101111" => data <= "000000";
				when "10111011110000" => data <= "000000";
				when "10111011110001" => data <= "000000";
				when "10111011110010" => data <= "000000";
				when "10111011110011" => data <= "000000";
				when "10111011110100" => data <= "000000";
				when "10111011110101" => data <= "000000";
				when "10111011110110" => data <= "000000";
				when "10111011110111" => data <= "000000";
				when "10111011111000" => data <= "000000";
				when "10111011111001" => data <= "000000";
				when "10111011111010" => data <= "000000";
				when "10111011111011" => data <= "000000";
				when "10111011111100" => data <= "000000";
				when "10111011111101" => data <= "000000";
				when "10111011111110" => data <= "000000";
				when "10111011111111" => data <= "000000";
				when "10111100000000" => data <= "000000";
				when "10111100000001" => data <= "000000";
				when "10111100000010" => data <= "000000";
				when "10111100000011" => data <= "000000";
				when "10111100000100" => data <= "000000";
				when "10111100000101" => data <= "000000";
				when "10111100000110" => data <= "000000";
				when "10111100000111" => data <= "000000";
				when "10111100001000" => data <= "000000";
				when "10111100001001" => data <= "000000";
				when "10111100001010" => data <= "000000";
				when "10111100001011" => data <= "000000";
				when "10111100001100" => data <= "000000";
				when "10111100001101" => data <= "000000";
				when "10111100001110" => data <= "000000";
				when "10111100001111" => data <= "000000";
				when "10111100010000" => data <= "000000";
				when "10111100010001" => data <= "000000";
				when "10111100010010" => data <= "000000";
				when "10111100010011" => data <= "000000";
				when "10111100010100" => data <= "000000";
				when "10111100010101" => data <= "000000";
				when "10111100010110" => data <= "000000";
				when "10111100010111" => data <= "000000";
				when "10111100011000" => data <= "000000";
				when "10111100011001" => data <= "000000";
				when "10111100011010" => data <= "000000";
				when "10111100011011" => data <= "000000";
				when "10111100011100" => data <= "000000";
				when "10111100011101" => data <= "000000";
				when "10111100011110" => data <= "000000";
				when "10111100011111" => data <= "000000";
				when "10111100100000" => data <= "000000";
				when "10111100100001" => data <= "000000";
				when "10111100100010" => data <= "000000";
				when "10111100100011" => data <= "000000";
				when "10111100100100" => data <= "000000";
				when "10111100100101" => data <= "000000";
				when "10111100100110" => data <= "000000";
				when "10111100100111" => data <= "000000";
				when "10111100101000" => data <= "000000";
				when "10111100101001" => data <= "000000";
				when "10111100101010" => data <= "000000";
				when "10111100101011" => data <= "000000";
				when "10111100101100" => data <= "000000";
				when "10111100101101" => data <= "000000";
				when "10111100101110" => data <= "000000";
				when "10111100101111" => data <= "000000";
				when "10111100110000" => data <= "000000";
				when "10111100110001" => data <= "000000";
				when "10111100110010" => data <= "000000";
				when "10111100110011" => data <= "000000";
				when "10111100110100" => data <= "000000";
				when "10111100110101" => data <= "000000";
				when "10111100110110" => data <= "000000";
				when "10111100110111" => data <= "000000";
				when "10111100111000" => data <= "000000";
				when "10111100111001" => data <= "000000";
				when "10111100111010" => data <= "000000";
				when "10111100111011" => data <= "000000";
				when "10111100111100" => data <= "000000";
				when "10111100111101" => data <= "000000";
				when "10111100111110" => data <= "000000";
				when "10111100111111" => data <= "000000";
				when "10111101000000" => data <= "000000";
				when "10111101000001" => data <= "000000";
				when "10111101000010" => data <= "000000";
				when "10111101000011" => data <= "000000";
				when "10111101000100" => data <= "000000";
				when "10111101000101" => data <= "000000";
				when "10111101000110" => data <= "000000";
				when "10111101000111" => data <= "000000";
				when "10111101001000" => data <= "000000";
				when "10111101001001" => data <= "000000";
				when "10111101001010" => data <= "000000";
				when "10111101001011" => data <= "000000";
				when "10111101001100" => data <= "000000";
				when "10111101001101" => data <= "000000";
				when "10111101001110" => data <= "000000";
				when "10111101001111" => data <= "000000";
				when "10111101010000" => data <= "000000";
				when "10111101010001" => data <= "000000";
				when "10111101010010" => data <= "000000";
				when "10111101010011" => data <= "000000";
				when "10111101010100" => data <= "000000";
				when "10111101010101" => data <= "000000";
				when "10111101010110" => data <= "000000";
				when "10111101010111" => data <= "000000";
				when "10111101011000" => data <= "000000";
				when "10111101011001" => data <= "000000";
				when "10111101011010" => data <= "000000";
				when "10111101011011" => data <= "000000";
				when "10111101011100" => data <= "000000";
				when "10111101011101" => data <= "000000";
				when "10111101011110" => data <= "000000";
				when "10111101011111" => data <= "000000";
				when "10111101100000" => data <= "000000";
				when "10111101100001" => data <= "000000";
				when "10111101100010" => data <= "000000";
				when "10111101100011" => data <= "000000";
				when "10111101100100" => data <= "000000";
				when "10111101100101" => data <= "000000";
				when "10111101100110" => data <= "000000";
				when "10111101100111" => data <= "000000";
				when "10111101101000" => data <= "000000";
				when "10111101101001" => data <= "000000";
				when "10111101101010" => data <= "000000";
				when "10111101101011" => data <= "000000";
				when "10111101101100" => data <= "000000";
				when "10111101101101" => data <= "000000";
				when "10111101101110" => data <= "000000";
				when "10111101101111" => data <= "000000";
				when "10111101110000" => data <= "000000";
				when "10111101110001" => data <= "000000";
				when "10111101110010" => data <= "000000";
				when "10111101110011" => data <= "000000";
				when "10111101110100" => data <= "000000";
				when "10111101110101" => data <= "000000";
				when "10111101110110" => data <= "000000";
				when "10111101110111" => data <= "000000";
				when "10111101111000" => data <= "000000";
				when "10111101111001" => data <= "000000";
				when "10111101111010" => data <= "000000";
				when "10111101111011" => data <= "000000";
				when "10111101111100" => data <= "000000";
				when "10111101111101" => data <= "000000";
				when "10111101111110" => data <= "000000";
				when "10111101111111" => data <= "000000";
				when "10111110000000" => data <= "000000";
				when "10111110000001" => data <= "000000";
				when "10111110000010" => data <= "000000";
				when "10111110000011" => data <= "000000";
				when "10111110000100" => data <= "000000";
				when "10111110000101" => data <= "000000";
				when "10111110000110" => data <= "000000";
				when "10111110000111" => data <= "000000";
				when "10111110001000" => data <= "000000";
				when "10111110001001" => data <= "000000";
				when "10111110001010" => data <= "000000";
				when "10111110001011" => data <= "000000";
				when "10111110001100" => data <= "000000";
				when "10111110001101" => data <= "000000";
				when "10111110001110" => data <= "000000";
				when "10111110001111" => data <= "000000";
				when "10111110010000" => data <= "000000";
				when "10111110010001" => data <= "000000";
				when "10111110010010" => data <= "000000";
				when "10111110010011" => data <= "000000";
				when "10111110010100" => data <= "000000";
				when "10111110010101" => data <= "000000";
				when "10111110010110" => data <= "000000";
				when "10111110010111" => data <= "000000";
				when "10111110011000" => data <= "000000";
				when "10111110011001" => data <= "000000";
				when "10111110011010" => data <= "000000";
				when "10111110011011" => data <= "000000";
				when "10111110011100" => data <= "000000";
				when "10111110011101" => data <= "000000";
				when "10111110011110" => data <= "000000";
				when "10111110011111" => data <= "000000";
				when "10111110100000" => data <= "000000";
				when "10111110100001" => data <= "000000";
				when "10111110100010" => data <= "000000";
				when "10111110100011" => data <= "000000";
				when "10111110100100" => data <= "000000";
				when "10111110100101" => data <= "000000";
				when "10111110100110" => data <= "000000";
				when "10111110100111" => data <= "000000";
				when "10111110101000" => data <= "000000";
				when "10111110101001" => data <= "000000";
				when "10111110101010" => data <= "000000";
				when "10111110101011" => data <= "000000";
				when "10111110101100" => data <= "000000";
				when "10111110101101" => data <= "000000";
				when "10111110101110" => data <= "000000";
				when "10111110101111" => data <= "000000";
				when "10111110110000" => data <= "000000";
				when "10111110110001" => data <= "000000";
				when "10111110110010" => data <= "000000";
				when "10111110110011" => data <= "000000";
				when "10111110110100" => data <= "000000";
				when "10111110110101" => data <= "000000";
				when "10111110110110" => data <= "000000";
				when "10111110110111" => data <= "000000";
				when "10111110111000" => data <= "000000";
				when "10111110111001" => data <= "000000";
				when "10111110111010" => data <= "000000";
				when "10111110111011" => data <= "000000";
				when "10111110111100" => data <= "000000";
				when "10111110111101" => data <= "000000";
				when "10111110111110" => data <= "000000";
				when "10111110111111" => data <= "000000";
				when "10111111000000" => data <= "000000";
				when "10111111000001" => data <= "000000";
				when "10111111000010" => data <= "000000";
				when "10111111000011" => data <= "000000";
				when "10111111000100" => data <= "000000";
				when "10111111000101" => data <= "000000";
				when "10111111000110" => data <= "000000";
				when "10111111000111" => data <= "000000";
				when "10111111001000" => data <= "000000";
				when "10111111001001" => data <= "000000";
				when "10111111001010" => data <= "000000";
				when "10111111001011" => data <= "000000";
				when "10111111001100" => data <= "000000";
				when "10111111001101" => data <= "000000";
				when "10111111001110" => data <= "000000";
				when "10111111001111" => data <= "000000";
				when "10111111010000" => data <= "000000";
				when "10111111010001" => data <= "000000";
				when "10111111010010" => data <= "000000";
				when "10111111010011" => data <= "000000";
				when "10111111010100" => data <= "000000";
				when "10111111010101" => data <= "000000";
				when "10111111010110" => data <= "000000";
				when "10111111010111" => data <= "000000";
				when "10111111011000" => data <= "000000";
				when "10111111011001" => data <= "000000";
				when "10111111011010" => data <= "000000";
				when "10111111011011" => data <= "000000";
				when "10111111011100" => data <= "000000";
				when "10111111011101" => data <= "000000";
				when "10111111011110" => data <= "000000";
				when "10111111011111" => data <= "000000";
				when "10111111100000" => data <= "000000";
				when "10111111100001" => data <= "000000";
				when "10111111100010" => data <= "000000";
				when "10111111100011" => data <= "000000";
				when "10111111100100" => data <= "000000";
				when "10111111100101" => data <= "000000";
				when "10111111100110" => data <= "000000";
				when "10111111100111" => data <= "000000";
				when "10111111101000" => data <= "000000";
				when "10111111101001" => data <= "000000";
				when "10111111101010" => data <= "000000";
				when "10111111101011" => data <= "000000";
				when "10111111101100" => data <= "000000";
				when "10111111101101" => data <= "000000";
				when "10111111101110" => data <= "000000";
				when "10111111101111" => data <= "000000";
				when "10111111110000" => data <= "000000";
				when "10111111110001" => data <= "000000";
				when "10111111110010" => data <= "000000";
				when "10111111110011" => data <= "000000";
				when "10111111110100" => data <= "000000";
				when "10111111110101" => data <= "000000";
				when "10111111110110" => data <= "000000";
				when "10111111110111" => data <= "000000";
				when "10111111111000" => data <= "000000";
				when "10111111111001" => data <= "000000";
				when "10111111111010" => data <= "000000";
				when "10111111111011" => data <= "000000";
				when "10111111111100" => data <= "000000";
				when "10111111111101" => data <= "000000";
				when "10111111111110" => data <= "000000";
				when "10111111111111" => data <= "000000";
				when others => data <= "000000";
			end case;
              		end if; 
              	end process; 
              end;