library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity rom is 
                 	port(
                		outglobal_o : in std_logic;
                		addr_x : in std_logic_vector(7 downto 0);
                		addr_y : in std_logic_vector(7 downto 0);
                		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
                	);
                end;

                architecture sim of rom is
                signal addr : std_logic_vector(15 downto 0);

                begin
                	addr (15 downto 8) <= addr_x;
                	addr (7 downto 0) <= addr_y;
                	process(outglobal_o) begin
                		if rising_edge(outglobal_o) then
                			case addr is
				when "0000111100101010" => data <= "111111";
				when "0000111100101011" => data <= "111111";
				when "0000111100101100" => data <= "111111";
				when "0000111100101101" => data <= "111111";
				when "0000111100101110" => data <= "111111";
				when "0000111100101111" => data <= "111111";
				when "0000111100110000" => data <= "111111";
				when "0000111100110001" => data <= "111111";
				when "0000111100111100" => data <= "111111";
				when "0000111100111101" => data <= "111111";
				when "0000111100111110" => data <= "111111";
				when "0000111100111111" => data <= "111111";
				when "0000111101000000" => data <= "111111";
				when "0000111101000001" => data <= "111111";
				when "0000111101000010" => data <= "111111";
				when "0000111101000011" => data <= "111111";
				when "0000111101000100" => data <= "111111";
				when "0000111101000101" => data <= "111111";
				when "0000111101001101" => data <= "111111";
				when "0000111101001110" => data <= "111111";
				when "0000111101001111" => data <= "111111";
				when "0000111101010000" => data <= "111111";
				when "0000111101010001" => data <= "111111";
				when "0000111101010010" => data <= "111111";
				when "0000111101010011" => data <= "111111";
				when "0000111101010100" => data <= "111111";
				when "0000111101010101" => data <= "111111";
				when "0000111101010110" => data <= "111111";
				when "0000111101010111" => data <= "111111";
				when "0000111101011000" => data <= "111111";
				when "0000111101100000" => data <= "111111";
				when "0000111101100001" => data <= "111111";
				when "0000111101100010" => data <= "111111";
				when "0000111101100011" => data <= "111111";
				when "0000111101100100" => data <= "111111";
				when "0000111101100101" => data <= "111111";
				when "0000111101100110" => data <= "111111";
				when "0000111101100111" => data <= "111111";
				when "0000111101110100" => data <= "111111";
				when "0000111101110101" => data <= "111111";
				when "0000111101110110" => data <= "111111";
				when "0000111101110111" => data <= "111111";
				when "0000111101111000" => data <= "111111";
				when "0000111101111001" => data <= "111111";
				when "0000111101111010" => data <= "111111";
				when "0000111101111011" => data <= "111111";
				when "0001000000101001" => data <= "111111";
				when "0001000000101010" => data <= "010010";
				when "0001000000101011" => data <= "010010";
				when "0001000000101100" => data <= "010010";
				when "0001000000101101" => data <= "010010";
				when "0001000000101110" => data <= "010010";
				when "0001000000101111" => data <= "010010";
				when "0001000000110000" => data <= "010010";
				when "0001000000110001" => data <= "010010";
				when "0001000000110010" => data <= "111111";
				when "0001000000111011" => data <= "111111";
				when "0001000000111100" => data <= "010010";
				when "0001000000111101" => data <= "010010";
				when "0001000000111110" => data <= "010010";
				when "0001000000111111" => data <= "010010";
				when "0001000001000000" => data <= "010010";
				when "0001000001000001" => data <= "010010";
				when "0001000001000010" => data <= "010010";
				when "0001000001000011" => data <= "010010";
				when "0001000001000100" => data <= "010010";
				when "0001000001000101" => data <= "010010";
				when "0001000001000110" => data <= "111111";
				when "0001000001001100" => data <= "111111";
				when "0001000001001101" => data <= "010010";
				when "0001000001001110" => data <= "010010";
				when "0001000001001111" => data <= "010010";
				when "0001000001010000" => data <= "010010";
				when "0001000001010001" => data <= "010010";
				when "0001000001010010" => data <= "010010";
				when "0001000001010011" => data <= "010010";
				when "0001000001010100" => data <= "010010";
				when "0001000001010101" => data <= "010010";
				when "0001000001010110" => data <= "010010";
				when "0001000001010111" => data <= "010010";
				when "0001000001011000" => data <= "010010";
				when "0001000001011001" => data <= "111111";
				when "0001000001011111" => data <= "111111";
				when "0001000001100000" => data <= "010010";
				when "0001000001100001" => data <= "010010";
				when "0001000001100010" => data <= "010010";
				when "0001000001100011" => data <= "010010";
				when "0001000001100100" => data <= "010010";
				when "0001000001100101" => data <= "010010";
				when "0001000001100110" => data <= "010010";
				when "0001000001100111" => data <= "010010";
				when "0001000001101000" => data <= "111111";
				when "0001000001110011" => data <= "111111";
				when "0001000001110100" => data <= "010010";
				when "0001000001110101" => data <= "010010";
				when "0001000001110110" => data <= "010010";
				when "0001000001110111" => data <= "010010";
				when "0001000001111000" => data <= "010010";
				when "0001000001111001" => data <= "010010";
				when "0001000001111010" => data <= "010010";
				when "0001000001111011" => data <= "010010";
				when "0001000001111100" => data <= "111111";
				when "0001000100101001" => data <= "111111";
				when "0001000100101010" => data <= "010010";
				when "0001000100101011" => data <= "010010";
				when "0001000100101100" => data <= "010010";
				when "0001000100101101" => data <= "010010";
				when "0001000100101110" => data <= "010010";
				when "0001000100101111" => data <= "010010";
				when "0001000100110000" => data <= "010010";
				when "0001000100110001" => data <= "010010";
				when "0001000100110010" => data <= "111111";
				when "0001000100110011" => data <= "111111";
				when "0001000100111011" => data <= "111111";
				when "0001000100111100" => data <= "010010";
				when "0001000100111101" => data <= "010010";
				when "0001000100111110" => data <= "010010";
				when "0001000100111111" => data <= "010010";
				when "0001000101000000" => data <= "010010";
				when "0001000101000001" => data <= "010010";
				when "0001000101000010" => data <= "010010";
				when "0001000101000011" => data <= "010010";
				when "0001000101000100" => data <= "010010";
				when "0001000101000101" => data <= "010010";
				when "0001000101000110" => data <= "111111";
				when "0001000101001100" => data <= "111111";
				when "0001000101001101" => data <= "010010";
				when "0001000101001110" => data <= "010010";
				when "0001000101001111" => data <= "010010";
				when "0001000101010000" => data <= "010010";
				when "0001000101010001" => data <= "010010";
				when "0001000101010010" => data <= "010010";
				when "0001000101010011" => data <= "010010";
				when "0001000101010100" => data <= "010010";
				when "0001000101010101" => data <= "010010";
				when "0001000101010110" => data <= "010010";
				when "0001000101010111" => data <= "010010";
				when "0001000101011000" => data <= "010010";
				when "0001000101011001" => data <= "111111";
				when "0001000101011111" => data <= "111111";
				when "0001000101100000" => data <= "010010";
				when "0001000101100001" => data <= "010010";
				when "0001000101100010" => data <= "010010";
				when "0001000101100011" => data <= "010010";
				when "0001000101100100" => data <= "010010";
				when "0001000101100101" => data <= "010010";
				when "0001000101100110" => data <= "010010";
				when "0001000101100111" => data <= "010010";
				when "0001000101101000" => data <= "111111";
				when "0001000101101001" => data <= "111111";
				when "0001000101110010" => data <= "111111";
				when "0001000101110011" => data <= "010010";
				when "0001000101110100" => data <= "010010";
				when "0001000101110101" => data <= "010010";
				when "0001000101110110" => data <= "010010";
				when "0001000101110111" => data <= "010010";
				when "0001000101111000" => data <= "010010";
				when "0001000101111001" => data <= "010010";
				when "0001000101111010" => data <= "010010";
				when "0001000101111011" => data <= "010010";
				when "0001000101111100" => data <= "010010";
				when "0001000101111101" => data <= "111111";
				when "0001001000101001" => data <= "111111";
				when "0001001000101010" => data <= "010010";
				when "0001001000101011" => data <= "010010";
				when "0001001000101100" => data <= "111111";
				when "0001001000101101" => data <= "111111";
				when "0001001000101110" => data <= "111111";
				when "0001001000101111" => data <= "111111";
				when "0001001000110000" => data <= "111111";
				when "0001001000110001" => data <= "111111";
				when "0001001000110010" => data <= "010010";
				when "0001001000110011" => data <= "010010";
				when "0001001000110100" => data <= "111111";
				when "0001001000111011" => data <= "111111";
				when "0001001000111100" => data <= "010010";
				when "0001001000111101" => data <= "010010";
				when "0001001000111110" => data <= "111111";
				when "0001001000111111" => data <= "111111";
				when "0001001001000000" => data <= "111111";
				when "0001001001000001" => data <= "111111";
				when "0001001001000010" => data <= "111111";
				when "0001001001000011" => data <= "111111";
				when "0001001001000100" => data <= "111111";
				when "0001001001000101" => data <= "111111";
				when "0001001001001101" => data <= "111111";
				when "0001001001001110" => data <= "111111";
				when "0001001001001111" => data <= "111111";
				when "0001001001010000" => data <= "111111";
				when "0001001001010001" => data <= "111111";
				when "0001001001010010" => data <= "010010";
				when "0001001001010011" => data <= "010010";
				when "0001001001010100" => data <= "111111";
				when "0001001001010101" => data <= "111111";
				when "0001001001010110" => data <= "111111";
				when "0001001001010111" => data <= "111111";
				when "0001001001011000" => data <= "111111";
				when "0001001001011111" => data <= "111111";
				when "0001001001100000" => data <= "010010";
				when "0001001001100001" => data <= "010010";
				when "0001001001100010" => data <= "111111";
				when "0001001001100011" => data <= "111111";
				when "0001001001100100" => data <= "111111";
				when "0001001001100101" => data <= "111111";
				when "0001001001100110" => data <= "111111";
				when "0001001001100111" => data <= "111111";
				when "0001001001101000" => data <= "010010";
				when "0001001001101001" => data <= "010010";
				when "0001001001101010" => data <= "111111";
				when "0001001001110001" => data <= "111111";
				when "0001001001110010" => data <= "010010";
				when "0001001001110011" => data <= "010010";
				when "0001001001110100" => data <= "111111";
				when "0001001001110101" => data <= "111111";
				when "0001001001110110" => data <= "111111";
				when "0001001001110111" => data <= "111111";
				when "0001001001111000" => data <= "111111";
				when "0001001001111001" => data <= "111111";
				when "0001001001111010" => data <= "111111";
				when "0001001001111011" => data <= "111111";
				when "0001001001111100" => data <= "010010";
				when "0001001001111101" => data <= "010010";
				when "0001001001111110" => data <= "111111";
				when "0001001100101001" => data <= "111111";
				when "0001001100101010" => data <= "010010";
				when "0001001100101011" => data <= "010010";
				when "0001001100101100" => data <= "111111";
				when "0001001100110001" => data <= "111111";
				when "0001001100110010" => data <= "010010";
				when "0001001100110011" => data <= "010010";
				when "0001001100110100" => data <= "111111";
				when "0001001100111011" => data <= "111111";
				when "0001001100111100" => data <= "010010";
				when "0001001100111101" => data <= "010010";
				when "0001001100111110" => data <= "111111";
				when "0001001101010001" => data <= "111111";
				when "0001001101010010" => data <= "010010";
				when "0001001101010011" => data <= "010010";
				when "0001001101010100" => data <= "111111";
				when "0001001101011111" => data <= "111111";
				when "0001001101100000" => data <= "010010";
				when "0001001101100001" => data <= "010010";
				when "0001001101100010" => data <= "111111";
				when "0001001101100111" => data <= "111111";
				when "0001001101101000" => data <= "010010";
				when "0001001101101001" => data <= "010010";
				when "0001001101101010" => data <= "111111";
				when "0001001101110001" => data <= "111111";
				when "0001001101110010" => data <= "010010";
				when "0001001101110011" => data <= "010010";
				when "0001001101110100" => data <= "111111";
				when "0001001101111011" => data <= "111111";
				when "0001001101111100" => data <= "010010";
				when "0001001101111101" => data <= "010010";
				when "0001001101111110" => data <= "111111";
				when "0001010000101001" => data <= "111111";
				when "0001010000101010" => data <= "010010";
				when "0001010000101011" => data <= "010010";
				when "0001010000101100" => data <= "111111";
				when "0001010000110001" => data <= "111111";
				when "0001010000110010" => data <= "010010";
				when "0001010000110011" => data <= "010010";
				when "0001010000110100" => data <= "111111";
				when "0001010000111011" => data <= "111111";
				when "0001010000111100" => data <= "010010";
				when "0001010000111101" => data <= "010010";
				when "0001010000111110" => data <= "111111";
				when "0001010001010001" => data <= "111111";
				when "0001010001010010" => data <= "010010";
				when "0001010001010011" => data <= "010010";
				when "0001010001010100" => data <= "111111";
				when "0001010001011111" => data <= "111111";
				when "0001010001100000" => data <= "010010";
				when "0001010001100001" => data <= "010010";
				when "0001010001100010" => data <= "111111";
				when "0001010001100111" => data <= "111111";
				when "0001010001101000" => data <= "010010";
				when "0001010001101001" => data <= "010010";
				when "0001010001101010" => data <= "111111";
				when "0001010001110001" => data <= "111111";
				when "0001010001110010" => data <= "010010";
				when "0001010001110011" => data <= "010010";
				when "0001010001110100" => data <= "111111";
				when "0001010001111011" => data <= "111111";
				when "0001010001111100" => data <= "010010";
				when "0001010001111101" => data <= "010010";
				when "0001010001111110" => data <= "111111";
				when "0001010100101001" => data <= "111111";
				when "0001010100101010" => data <= "100010";
				when "0001010100101011" => data <= "100010";
				when "0001010100101100" => data <= "111111";
				when "0001010100110001" => data <= "111111";
				when "0001010100110010" => data <= "100010";
				when "0001010100110011" => data <= "100010";
				when "0001010100110100" => data <= "111111";
				when "0001010100111011" => data <= "111111";
				when "0001010100111100" => data <= "100010";
				when "0001010100111101" => data <= "100010";
				when "0001010100111110" => data <= "111111";
				when "0001010101010001" => data <= "111111";
				when "0001010101010010" => data <= "100010";
				when "0001010101010011" => data <= "100010";
				when "0001010101010100" => data <= "111111";
				when "0001010101011111" => data <= "111111";
				when "0001010101100000" => data <= "100010";
				when "0001010101100001" => data <= "100010";
				when "0001010101100010" => data <= "111111";
				when "0001010101100111" => data <= "111111";
				when "0001010101101000" => data <= "100010";
				when "0001010101101001" => data <= "100010";
				when "0001010101101010" => data <= "111111";
				when "0001010101110001" => data <= "111111";
				when "0001010101110010" => data <= "100010";
				when "0001010101110011" => data <= "100010";
				when "0001010101110100" => data <= "111111";
				when "0001010101111011" => data <= "111111";
				when "0001010101111100" => data <= "100010";
				when "0001010101111101" => data <= "100010";
				when "0001010101111110" => data <= "111111";
				when "0001011000101001" => data <= "111111";
				when "0001011000101010" => data <= "100010";
				when "0001011000101011" => data <= "100010";
				when "0001011000101100" => data <= "111111";
				when "0001011000110001" => data <= "111111";
				when "0001011000110010" => data <= "100010";
				when "0001011000110011" => data <= "100010";
				when "0001011000110100" => data <= "111111";
				when "0001011000111011" => data <= "111111";
				when "0001011000111100" => data <= "100010";
				when "0001011000111101" => data <= "100010";
				when "0001011000111110" => data <= "111111";
				when "0001011001010001" => data <= "111111";
				when "0001011001010010" => data <= "100010";
				when "0001011001010011" => data <= "100010";
				when "0001011001010100" => data <= "111111";
				when "0001011001011111" => data <= "111111";
				when "0001011001100000" => data <= "100010";
				when "0001011001100001" => data <= "100010";
				when "0001011001100010" => data <= "111111";
				when "0001011001100111" => data <= "111111";
				when "0001011001101000" => data <= "100010";
				when "0001011001101001" => data <= "100010";
				when "0001011001101010" => data <= "111111";
				when "0001011001110001" => data <= "111111";
				when "0001011001110010" => data <= "100010";
				when "0001011001110011" => data <= "100010";
				when "0001011001110100" => data <= "111111";
				when "0001011001111011" => data <= "111111";
				when "0001011001111100" => data <= "100010";
				when "0001011001111101" => data <= "100010";
				when "0001011001111110" => data <= "111111";
				when "0001011100101001" => data <= "111111";
				when "0001011100101010" => data <= "100010";
				when "0001011100101011" => data <= "100010";
				when "0001011100101100" => data <= "111111";
				when "0001011100101101" => data <= "111111";
				when "0001011100101110" => data <= "111111";
				when "0001011100101111" => data <= "111111";
				when "0001011100110000" => data <= "111111";
				when "0001011100110001" => data <= "111111";
				when "0001011100110010" => data <= "100010";
				when "0001011100110011" => data <= "100010";
				when "0001011100110100" => data <= "111111";
				when "0001011100111011" => data <= "111111";
				when "0001011100111100" => data <= "100010";
				when "0001011100111101" => data <= "100010";
				when "0001011100111110" => data <= "111111";
				when "0001011100111111" => data <= "111111";
				when "0001011101000000" => data <= "111111";
				when "0001011101000001" => data <= "111111";
				when "0001011101000010" => data <= "111111";
				when "0001011101000011" => data <= "111111";
				when "0001011101010001" => data <= "111111";
				when "0001011101010010" => data <= "100010";
				when "0001011101010011" => data <= "100010";
				when "0001011101010100" => data <= "111111";
				when "0001011101011111" => data <= "111111";
				when "0001011101100000" => data <= "100010";
				when "0001011101100001" => data <= "100010";
				when "0001011101100010" => data <= "111111";
				when "0001011101100011" => data <= "111111";
				when "0001011101100100" => data <= "111111";
				when "0001011101100101" => data <= "111111";
				when "0001011101100110" => data <= "111111";
				when "0001011101100111" => data <= "111111";
				when "0001011101101000" => data <= "100010";
				when "0001011101101001" => data <= "100010";
				when "0001011101101010" => data <= "111111";
				when "0001011101110001" => data <= "111111";
				when "0001011101110010" => data <= "100010";
				when "0001011101110011" => data <= "100010";
				when "0001011101110100" => data <= "111111";
				when "0001011101111011" => data <= "111111";
				when "0001011101111100" => data <= "100010";
				when "0001011101111101" => data <= "100010";
				when "0001011101111110" => data <= "111111";
				when "0001100000101001" => data <= "111111";
				when "0001100000101010" => data <= "100010";
				when "0001100000101011" => data <= "100010";
				when "0001100000101100" => data <= "100010";
				when "0001100000101101" => data <= "100010";
				when "0001100000101110" => data <= "100010";
				when "0001100000101111" => data <= "100010";
				when "0001100000110000" => data <= "100010";
				when "0001100000110001" => data <= "100010";
				when "0001100000110010" => data <= "111111";
				when "0001100000110011" => data <= "111111";
				when "0001100000111011" => data <= "111111";
				when "0001100000111100" => data <= "100010";
				when "0001100000111101" => data <= "100010";
				when "0001100000111110" => data <= "100010";
				when "0001100000111111" => data <= "100010";
				when "0001100001000000" => data <= "100010";
				when "0001100001000001" => data <= "100010";
				when "0001100001000010" => data <= "100010";
				when "0001100001000011" => data <= "100010";
				when "0001100001000100" => data <= "111111";
				when "0001100001010001" => data <= "111111";
				when "0001100001010010" => data <= "100010";
				when "0001100001010011" => data <= "100010";
				when "0001100001010100" => data <= "111111";
				when "0001100001011111" => data <= "111111";
				when "0001100001100000" => data <= "100010";
				when "0001100001100001" => data <= "100010";
				when "0001100001100010" => data <= "100010";
				when "0001100001100011" => data <= "100010";
				when "0001100001100100" => data <= "100010";
				when "0001100001100101" => data <= "100010";
				when "0001100001100110" => data <= "100010";
				when "0001100001100111" => data <= "100010";
				when "0001100001101000" => data <= "111111";
				when "0001100001101001" => data <= "111111";
				when "0001100001110001" => data <= "111111";
				when "0001100001110010" => data <= "100010";
				when "0001100001110011" => data <= "100010";
				when "0001100001110100" => data <= "111111";
				when "0001100001111011" => data <= "111111";
				when "0001100001111100" => data <= "100010";
				when "0001100001111101" => data <= "100010";
				when "0001100001111110" => data <= "111111";
				when "0001100100101001" => data <= "111111";
				when "0001100100101010" => data <= "100010";
				when "0001100100101011" => data <= "100010";
				when "0001100100101100" => data <= "100010";
				when "0001100100101101" => data <= "100010";
				when "0001100100101110" => data <= "100010";
				when "0001100100101111" => data <= "100010";
				when "0001100100110000" => data <= "100010";
				when "0001100100110001" => data <= "100010";
				when "0001100100110010" => data <= "111111";
				when "0001100100111011" => data <= "111111";
				when "0001100100111100" => data <= "100010";
				when "0001100100111101" => data <= "100010";
				when "0001100100111110" => data <= "100010";
				when "0001100100111111" => data <= "100010";
				when "0001100101000000" => data <= "100010";
				when "0001100101000001" => data <= "100010";
				when "0001100101000010" => data <= "100010";
				when "0001100101000011" => data <= "100010";
				when "0001100101000100" => data <= "111111";
				when "0001100101010001" => data <= "111111";
				when "0001100101010010" => data <= "100010";
				when "0001100101010011" => data <= "100010";
				when "0001100101010100" => data <= "111111";
				when "0001100101011111" => data <= "111111";
				when "0001100101100000" => data <= "100010";
				when "0001100101100001" => data <= "100010";
				when "0001100101100010" => data <= "100010";
				when "0001100101100011" => data <= "100010";
				when "0001100101100100" => data <= "100010";
				when "0001100101100101" => data <= "100010";
				when "0001100101100110" => data <= "100010";
				when "0001100101100111" => data <= "100010";
				when "0001100101101000" => data <= "111111";
				when "0001100101110001" => data <= "111111";
				when "0001100101110010" => data <= "100010";
				when "0001100101110011" => data <= "100010";
				when "0001100101110100" => data <= "111111";
				when "0001100101111011" => data <= "111111";
				when "0001100101111100" => data <= "100010";
				when "0001100101111101" => data <= "100010";
				when "0001100101111110" => data <= "111111";
				when "0001101000101001" => data <= "111111";
				when "0001101000101010" => data <= "100010";
				when "0001101000101011" => data <= "100010";
				when "0001101000101100" => data <= "111111";
				when "0001101000101101" => data <= "111111";
				when "0001101000101110" => data <= "111111";
				when "0001101000101111" => data <= "111111";
				when "0001101000110000" => data <= "111111";
				when "0001101000110001" => data <= "111111";
				when "0001101000110010" => data <= "100010";
				when "0001101000110011" => data <= "111111";
				when "0001101000111011" => data <= "111111";
				when "0001101000111100" => data <= "100010";
				when "0001101000111101" => data <= "100010";
				when "0001101000111110" => data <= "111111";
				when "0001101000111111" => data <= "111111";
				when "0001101001000000" => data <= "111111";
				when "0001101001000001" => data <= "111111";
				when "0001101001000010" => data <= "111111";
				when "0001101001000011" => data <= "111111";
				when "0001101001010001" => data <= "111111";
				when "0001101001010010" => data <= "100010";
				when "0001101001010011" => data <= "100010";
				when "0001101001010100" => data <= "111111";
				when "0001101001011111" => data <= "111111";
				when "0001101001100000" => data <= "100010";
				when "0001101001100001" => data <= "100010";
				when "0001101001100010" => data <= "111111";
				when "0001101001100011" => data <= "111111";
				when "0001101001100100" => data <= "111111";
				when "0001101001100101" => data <= "111111";
				when "0001101001100110" => data <= "111111";
				when "0001101001100111" => data <= "111111";
				when "0001101001101000" => data <= "100010";
				when "0001101001101001" => data <= "111111";
				when "0001101001110001" => data <= "111111";
				when "0001101001110010" => data <= "100010";
				when "0001101001110011" => data <= "100010";
				when "0001101001110100" => data <= "111111";
				when "0001101001111011" => data <= "111111";
				when "0001101001111100" => data <= "100010";
				when "0001101001111101" => data <= "100010";
				when "0001101001111110" => data <= "111111";
				when "0001101100101001" => data <= "111111";
				when "0001101100101010" => data <= "100010";
				when "0001101100101011" => data <= "100010";
				when "0001101100101100" => data <= "111111";
				when "0001101100110001" => data <= "111111";
				when "0001101100110010" => data <= "100010";
				when "0001101100110011" => data <= "100010";
				when "0001101100110100" => data <= "111111";
				when "0001101100111011" => data <= "111111";
				when "0001101100111100" => data <= "100010";
				when "0001101100111101" => data <= "100010";
				when "0001101100111110" => data <= "111111";
				when "0001101101010001" => data <= "111111";
				when "0001101101010010" => data <= "100010";
				when "0001101101010011" => data <= "100010";
				when "0001101101010100" => data <= "111111";
				when "0001101101011111" => data <= "111111";
				when "0001101101100000" => data <= "100010";
				when "0001101101100001" => data <= "100010";
				when "0001101101100010" => data <= "111111";
				when "0001101101100111" => data <= "111111";
				when "0001101101101000" => data <= "100010";
				when "0001101101101001" => data <= "100010";
				when "0001101101101010" => data <= "111111";
				when "0001101101110001" => data <= "111111";
				when "0001101101110010" => data <= "100010";
				when "0001101101110011" => data <= "100010";
				when "0001101101110100" => data <= "111111";
				when "0001101101111011" => data <= "111111";
				when "0001101101111100" => data <= "100010";
				when "0001101101111101" => data <= "100010";
				when "0001101101111110" => data <= "111111";
				when "0001110000101001" => data <= "111111";
				when "0001110000101010" => data <= "100010";
				when "0001110000101011" => data <= "100010";
				when "0001110000101100" => data <= "111111";
				when "0001110000110001" => data <= "111111";
				when "0001110000110010" => data <= "100010";
				when "0001110000110011" => data <= "100010";
				when "0001110000110100" => data <= "111111";
				when "0001110000111011" => data <= "111111";
				when "0001110000111100" => data <= "100010";
				when "0001110000111101" => data <= "100010";
				when "0001110000111110" => data <= "111111";
				when "0001110001010001" => data <= "111111";
				when "0001110001010010" => data <= "100010";
				when "0001110001010011" => data <= "100010";
				when "0001110001010100" => data <= "111111";
				when "0001110001011111" => data <= "111111";
				when "0001110001100000" => data <= "100010";
				when "0001110001100001" => data <= "100010";
				when "0001110001100010" => data <= "111111";
				when "0001110001100111" => data <= "111111";
				when "0001110001101000" => data <= "100010";
				when "0001110001101001" => data <= "100010";
				when "0001110001101010" => data <= "111111";
				when "0001110001110001" => data <= "111111";
				when "0001110001110010" => data <= "100010";
				when "0001110001110011" => data <= "100010";
				when "0001110001110100" => data <= "111111";
				when "0001110001111011" => data <= "111111";
				when "0001110001111100" => data <= "100010";
				when "0001110001111101" => data <= "100010";
				when "0001110001111110" => data <= "111111";
				when "0001110100101001" => data <= "111111";
				when "0001110100101010" => data <= "100010";
				when "0001110100101011" => data <= "100010";
				when "0001110100101100" => data <= "111111";
				when "0001110100110001" => data <= "111111";
				when "0001110100110010" => data <= "100010";
				when "0001110100110011" => data <= "100010";
				when "0001110100110100" => data <= "111111";
				when "0001110100111011" => data <= "111111";
				when "0001110100111100" => data <= "100010";
				when "0001110100111101" => data <= "100010";
				when "0001110100111110" => data <= "111111";
				when "0001110101010001" => data <= "111111";
				when "0001110101010010" => data <= "110010";
				when "0001110101010011" => data <= "110010";
				when "0001110101010100" => data <= "111111";
				when "0001110101011111" => data <= "111111";
				when "0001110101100000" => data <= "110010";
				when "0001110101100001" => data <= "110010";
				when "0001110101100010" => data <= "111111";
				when "0001110101100111" => data <= "111111";
				when "0001110101101000" => data <= "110010";
				when "0001110101101001" => data <= "110010";
				when "0001110101101010" => data <= "111111";
				when "0001110101110001" => data <= "111111";
				when "0001110101110010" => data <= "110010";
				when "0001110101110011" => data <= "110010";
				when "0001110101110100" => data <= "111111";
				when "0001110101111011" => data <= "111111";
				when "0001110101111100" => data <= "110010";
				when "0001110101111101" => data <= "110010";
				when "0001110101111110" => data <= "111111";
				when "0001111000101001" => data <= "111111";
				when "0001111000101010" => data <= "110010";
				when "0001111000101011" => data <= "110010";
				when "0001111000101100" => data <= "111111";
				when "0001111000110001" => data <= "111111";
				when "0001111000110010" => data <= "110010";
				when "0001111000110011" => data <= "110010";
				when "0001111000110100" => data <= "111111";
				when "0001111000111011" => data <= "111111";
				when "0001111000111100" => data <= "110010";
				when "0001111000111101" => data <= "110010";
				when "0001111000111110" => data <= "111111";
				when "0001111000111111" => data <= "111111";
				when "0001111001000000" => data <= "111111";
				when "0001111001000001" => data <= "111111";
				when "0001111001000010" => data <= "111111";
				when "0001111001000011" => data <= "111111";
				when "0001111001000100" => data <= "111111";
				when "0001111001000101" => data <= "111111";
				when "0001111001010001" => data <= "111111";
				when "0001111001010010" => data <= "110010";
				when "0001111001010011" => data <= "110010";
				when "0001111001010100" => data <= "111111";
				when "0001111001011111" => data <= "111111";
				when "0001111001100000" => data <= "110010";
				when "0001111001100001" => data <= "110010";
				when "0001111001100010" => data <= "111111";
				when "0001111001100111" => data <= "111111";
				when "0001111001101000" => data <= "110010";
				when "0001111001101001" => data <= "110010";
				when "0001111001101010" => data <= "111111";
				when "0001111001110001" => data <= "111111";
				when "0001111001110010" => data <= "110010";
				when "0001111001110011" => data <= "110010";
				when "0001111001110100" => data <= "111111";
				when "0001111001110101" => data <= "111111";
				when "0001111001110110" => data <= "111111";
				when "0001111001110111" => data <= "111111";
				when "0001111001111000" => data <= "111111";
				when "0001111001111001" => data <= "111111";
				when "0001111001111010" => data <= "111111";
				when "0001111001111011" => data <= "111111";
				when "0001111001111100" => data <= "110010";
				when "0001111001111101" => data <= "110010";
				when "0001111001111110" => data <= "111111";
				when "0001111100101001" => data <= "111111";
				when "0001111100101010" => data <= "110010";
				when "0001111100101011" => data <= "110010";
				when "0001111100101100" => data <= "111111";
				when "0001111100110001" => data <= "111111";
				when "0001111100110010" => data <= "110010";
				when "0001111100110011" => data <= "110010";
				when "0001111100110100" => data <= "111111";
				when "0001111100111011" => data <= "111111";
				when "0001111100111100" => data <= "110010";
				when "0001111100111101" => data <= "110010";
				when "0001111100111110" => data <= "110010";
				when "0001111100111111" => data <= "110010";
				when "0001111101000000" => data <= "110010";
				when "0001111101000001" => data <= "110010";
				when "0001111101000010" => data <= "110010";
				when "0001111101000011" => data <= "110010";
				when "0001111101000100" => data <= "110010";
				when "0001111101000101" => data <= "110010";
				when "0001111101000110" => data <= "111111";
				when "0001111101010001" => data <= "111111";
				when "0001111101010010" => data <= "110010";
				when "0001111101010011" => data <= "110010";
				when "0001111101010100" => data <= "111111";
				when "0001111101011111" => data <= "111111";
				when "0001111101100000" => data <= "110010";
				when "0001111101100001" => data <= "110010";
				when "0001111101100010" => data <= "111111";
				when "0001111101100111" => data <= "111111";
				when "0001111101101000" => data <= "110010";
				when "0001111101101001" => data <= "110010";
				when "0001111101101010" => data <= "111111";
				when "0001111101110010" => data <= "111111";
				when "0001111101110011" => data <= "110010";
				when "0001111101110100" => data <= "110010";
				when "0001111101110101" => data <= "110010";
				when "0001111101110110" => data <= "110010";
				when "0001111101110111" => data <= "110010";
				when "0001111101111000" => data <= "110010";
				when "0001111101111001" => data <= "110010";
				when "0001111101111010" => data <= "110010";
				when "0001111101111011" => data <= "110010";
				when "0001111101111100" => data <= "110010";
				when "0001111101111101" => data <= "111111";
				when "0010000000101001" => data <= "111111";
				when "0010000000101010" => data <= "110010";
				when "0010000000101011" => data <= "110010";
				when "0010000000101100" => data <= "111111";
				when "0010000000110001" => data <= "111111";
				when "0010000000110010" => data <= "110010";
				when "0010000000110011" => data <= "110010";
				when "0010000000110100" => data <= "111111";
				when "0010000000111011" => data <= "111111";
				when "0010000000111100" => data <= "110010";
				when "0010000000111101" => data <= "110010";
				when "0010000000111110" => data <= "110010";
				when "0010000000111111" => data <= "110010";
				when "0010000001000000" => data <= "110010";
				when "0010000001000001" => data <= "110010";
				when "0010000001000010" => data <= "110010";
				when "0010000001000011" => data <= "110010";
				when "0010000001000100" => data <= "110010";
				when "0010000001000101" => data <= "110010";
				when "0010000001000110" => data <= "111111";
				when "0010000001010001" => data <= "111111";
				when "0010000001010010" => data <= "110010";
				when "0010000001010011" => data <= "110010";
				when "0010000001010100" => data <= "111111";
				when "0010000001011111" => data <= "111111";
				when "0010000001100000" => data <= "110010";
				when "0010000001100001" => data <= "110010";
				when "0010000001100010" => data <= "111111";
				when "0010000001100111" => data <= "111111";
				when "0010000001101000" => data <= "110010";
				when "0010000001101001" => data <= "110010";
				when "0010000001101010" => data <= "111111";
				when "0010000001110011" => data <= "111111";
				when "0010000001110100" => data <= "110010";
				when "0010000001110101" => data <= "110010";
				when "0010000001110110" => data <= "110010";
				when "0010000001110111" => data <= "110010";
				when "0010000001111000" => data <= "110010";
				when "0010000001111001" => data <= "110010";
				when "0010000001111010" => data <= "110010";
				when "0010000001111011" => data <= "110010";
				when "0010000001111100" => data <= "111111";
				when "0010000100101010" => data <= "111111";
				when "0010000100101011" => data <= "111111";
				when "0010000100110010" => data <= "111111";
				when "0010000100110011" => data <= "111111";
				when "0010000100111100" => data <= "111111";
				when "0010000100111101" => data <= "111111";
				when "0010000100111110" => data <= "111111";
				when "0010000100111111" => data <= "111111";
				when "0010000101000000" => data <= "111111";
				when "0010000101000001" => data <= "111111";
				when "0010000101000010" => data <= "111111";
				when "0010000101000011" => data <= "111111";
				when "0010000101000100" => data <= "111111";
				when "0010000101000101" => data <= "111111";
				when "0010000101010010" => data <= "111111";
				when "0010000101010011" => data <= "111111";
				when "0010000101100000" => data <= "111111";
				when "0010000101100001" => data <= "111111";
				when "0010000101101000" => data <= "111111";
				when "0010000101101001" => data <= "111111";
				when "0010000101110100" => data <= "111111";
				when "0010000101110101" => data <= "111111";
				when "0010000101110110" => data <= "111111";
				when "0010000101110111" => data <= "111111";
				when "0010000101111000" => data <= "111111";
				when "0010000101111001" => data <= "111111";
				when "0010000101111010" => data <= "111111";
				when "0010000101111011" => data <= "111111";
				when "0010011000011100" => data <= "111111";
				when "0010011000011101" => data <= "111111";
				when "0010011000011110" => data <= "111111";
				when "0010011000011111" => data <= "111111";
				when "0010011000100000" => data <= "111111";
				when "0010011000100001" => data <= "111111";
				when "0010011000100010" => data <= "111111";
				when "0010011000100011" => data <= "111111";
				when "0010011000101100" => data <= "111111";
				when "0010011000101101" => data <= "111111";
				when "0010011000110100" => data <= "111111";
				when "0010011000110101" => data <= "111111";
				when "0010011000111100" => data <= "111111";
				when "0010011000111101" => data <= "111111";
				when "0010011001000100" => data <= "111111";
				when "0010011001000101" => data <= "111111";
				when "0010011001001011" => data <= "111111";
				when "0010011001001100" => data <= "111111";
				when "0010011001001101" => data <= "111111";
				when "0010011001001110" => data <= "111111";
				when "0010011001001111" => data <= "111111";
				when "0010011001010000" => data <= "111111";
				when "0010011001010001" => data <= "111111";
				when "0010011001010010" => data <= "111111";
				when "0010011001010011" => data <= "111111";
				when "0010011001010100" => data <= "111111";
				when "0010011001010101" => data <= "111111";
				when "0010011001010110" => data <= "111111";
				when "0010011001011101" => data <= "111111";
				when "0010011001011110" => data <= "111111";
				when "0010011001100101" => data <= "111111";
				when "0010011001100110" => data <= "111111";
				when "0010011001101101" => data <= "111111";
				when "0010011001101110" => data <= "111111";
				when "0010011001110101" => data <= "111111";
				when "0010011001110110" => data <= "111111";
				when "0010011001111110" => data <= "111111";
				when "0010011001111111" => data <= "111111";
				when "0010011010000110" => data <= "111111";
				when "0010011010000111" => data <= "111111";
				when "0010011100011011" => data <= "111111";
				when "0010011100011100" => data <= "010010";
				when "0010011100011101" => data <= "010010";
				when "0010011100011110" => data <= "010010";
				when "0010011100011111" => data <= "010010";
				when "0010011100100000" => data <= "010010";
				when "0010011100100001" => data <= "010010";
				when "0010011100100010" => data <= "010010";
				when "0010011100100011" => data <= "010010";
				when "0010011100100100" => data <= "111111";
				when "0010011100101011" => data <= "111111";
				when "0010011100101100" => data <= "010010";
				when "0010011100101101" => data <= "010010";
				when "0010011100101110" => data <= "111111";
				when "0010011100110011" => data <= "111111";
				when "0010011100110100" => data <= "010010";
				when "0010011100110101" => data <= "010010";
				when "0010011100110110" => data <= "111111";
				when "0010011100111011" => data <= "111111";
				when "0010011100111100" => data <= "010010";
				when "0010011100111101" => data <= "010010";
				when "0010011100111110" => data <= "111111";
				when "0010011101000011" => data <= "111111";
				when "0010011101000100" => data <= "010010";
				when "0010011101000101" => data <= "010010";
				when "0010011101000110" => data <= "111111";
				when "0010011101001010" => data <= "111111";
				when "0010011101001011" => data <= "010010";
				when "0010011101001100" => data <= "010010";
				when "0010011101001101" => data <= "010010";
				when "0010011101001110" => data <= "010010";
				when "0010011101001111" => data <= "010010";
				when "0010011101010000" => data <= "010010";
				when "0010011101010001" => data <= "010010";
				when "0010011101010010" => data <= "010010";
				when "0010011101010011" => data <= "010010";
				when "0010011101010100" => data <= "010010";
				when "0010011101010101" => data <= "010010";
				when "0010011101010110" => data <= "010010";
				when "0010011101010111" => data <= "111111";
				when "0010011101011100" => data <= "111111";
				when "0010011101011101" => data <= "010010";
				when "0010011101011110" => data <= "010010";
				when "0010011101011111" => data <= "111111";
				when "0010011101100100" => data <= "111111";
				when "0010011101100101" => data <= "010010";
				when "0010011101100110" => data <= "010010";
				when "0010011101100111" => data <= "111111";
				when "0010011101101100" => data <= "111111";
				when "0010011101101101" => data <= "010010";
				when "0010011101101110" => data <= "010010";
				when "0010011101101111" => data <= "111111";
				when "0010011101110100" => data <= "111111";
				when "0010011101110101" => data <= "010010";
				when "0010011101110110" => data <= "010010";
				when "0010011101110111" => data <= "111111";
				when "0010011101111101" => data <= "111111";
				when "0010011101111110" => data <= "010010";
				when "0010011101111111" => data <= "010010";
				when "0010011110000000" => data <= "111111";
				when "0010011110000101" => data <= "111111";
				when "0010011110000110" => data <= "010010";
				when "0010011110000111" => data <= "010010";
				when "0010011110001000" => data <= "111111";
				when "0010100000011011" => data <= "111111";
				when "0010100000011100" => data <= "010010";
				when "0010100000011101" => data <= "010010";
				when "0010100000011110" => data <= "010010";
				when "0010100000011111" => data <= "010010";
				when "0010100000100000" => data <= "010010";
				when "0010100000100001" => data <= "010010";
				when "0010100000100010" => data <= "010010";
				when "0010100000100011" => data <= "010010";
				when "0010100000100100" => data <= "111111";
				when "0010100000100101" => data <= "111111";
				when "0010100000101011" => data <= "111111";
				when "0010100000101100" => data <= "010010";
				when "0010100000101101" => data <= "010010";
				when "0010100000101110" => data <= "111111";
				when "0010100000110011" => data <= "111111";
				when "0010100000110100" => data <= "010010";
				when "0010100000110101" => data <= "010010";
				when "0010100000110110" => data <= "111111";
				when "0010100000111011" => data <= "111111";
				when "0010100000111100" => data <= "010010";
				when "0010100000111101" => data <= "010010";
				when "0010100000111110" => data <= "111111";
				when "0010100001000011" => data <= "111111";
				when "0010100001000100" => data <= "010010";
				when "0010100001000101" => data <= "010010";
				when "0010100001000110" => data <= "111111";
				when "0010100001001010" => data <= "111111";
				when "0010100001001011" => data <= "010010";
				when "0010100001001100" => data <= "010010";
				when "0010100001001101" => data <= "010010";
				when "0010100001001110" => data <= "010010";
				when "0010100001001111" => data <= "010010";
				when "0010100001010000" => data <= "010010";
				when "0010100001010001" => data <= "010010";
				when "0010100001010010" => data <= "010010";
				when "0010100001010011" => data <= "010010";
				when "0010100001010100" => data <= "010010";
				when "0010100001010101" => data <= "010010";
				when "0010100001010110" => data <= "010010";
				when "0010100001010111" => data <= "111111";
				when "0010100001011100" => data <= "111111";
				when "0010100001011101" => data <= "010010";
				when "0010100001011110" => data <= "010010";
				when "0010100001011111" => data <= "111111";
				when "0010100001100100" => data <= "111111";
				when "0010100001100101" => data <= "010010";
				when "0010100001100110" => data <= "010010";
				when "0010100001100111" => data <= "111111";
				when "0010100001101100" => data <= "111111";
				when "0010100001101101" => data <= "010010";
				when "0010100001101110" => data <= "010010";
				when "0010100001101111" => data <= "111111";
				when "0010100001110100" => data <= "111111";
				when "0010100001110101" => data <= "010010";
				when "0010100001110110" => data <= "010010";
				when "0010100001110111" => data <= "111111";
				when "0010100001111101" => data <= "111111";
				when "0010100001111110" => data <= "010010";
				when "0010100001111111" => data <= "010010";
				when "0010100010000000" => data <= "010010";
				when "0010100010000001" => data <= "111111";
				when "0010100010000100" => data <= "111111";
				when "0010100010000101" => data <= "010010";
				when "0010100010000110" => data <= "010010";
				when "0010100010000111" => data <= "010010";
				when "0010100010001000" => data <= "111111";
				when "0010100100011011" => data <= "111111";
				when "0010100100011100" => data <= "010010";
				when "0010100100011101" => data <= "010010";
				when "0010100100011110" => data <= "111111";
				when "0010100100011111" => data <= "111111";
				when "0010100100100000" => data <= "111111";
				when "0010100100100001" => data <= "111111";
				when "0010100100100010" => data <= "111111";
				when "0010100100100011" => data <= "111111";
				when "0010100100100100" => data <= "010010";
				when "0010100100100101" => data <= "010010";
				when "0010100100100110" => data <= "111111";
				when "0010100100101011" => data <= "111111";
				when "0010100100101100" => data <= "010010";
				when "0010100100101101" => data <= "010010";
				when "0010100100101110" => data <= "111111";
				when "0010100100110011" => data <= "111111";
				when "0010100100110100" => data <= "010010";
				when "0010100100110101" => data <= "010010";
				when "0010100100110110" => data <= "111111";
				when "0010100100111011" => data <= "111111";
				when "0010100100111100" => data <= "010010";
				when "0010100100111101" => data <= "010010";
				when "0010100100111110" => data <= "111111";
				when "0010100101000011" => data <= "111111";
				when "0010100101000100" => data <= "010010";
				when "0010100101000101" => data <= "010010";
				when "0010100101000110" => data <= "111111";
				when "0010100101001011" => data <= "111111";
				when "0010100101001100" => data <= "111111";
				when "0010100101001101" => data <= "111111";
				when "0010100101001110" => data <= "111111";
				when "0010100101001111" => data <= "111111";
				when "0010100101010000" => data <= "010010";
				when "0010100101010001" => data <= "010010";
				when "0010100101010010" => data <= "111111";
				when "0010100101010011" => data <= "111111";
				when "0010100101010100" => data <= "111111";
				when "0010100101010101" => data <= "111111";
				when "0010100101010110" => data <= "111111";
				when "0010100101011100" => data <= "111111";
				when "0010100101011101" => data <= "010010";
				when "0010100101011110" => data <= "010010";
				when "0010100101011111" => data <= "111111";
				when "0010100101100100" => data <= "111111";
				when "0010100101100101" => data <= "010010";
				when "0010100101100110" => data <= "010010";
				when "0010100101100111" => data <= "111111";
				when "0010100101101100" => data <= "111111";
				when "0010100101101101" => data <= "010010";
				when "0010100101101110" => data <= "010010";
				when "0010100101101111" => data <= "111111";
				when "0010100101110100" => data <= "111111";
				when "0010100101110101" => data <= "010010";
				when "0010100101110110" => data <= "010010";
				when "0010100101110111" => data <= "111111";
				when "0010100101111101" => data <= "111111";
				when "0010100101111110" => data <= "010010";
				when "0010100101111111" => data <= "010010";
				when "0010100110000000" => data <= "010010";
				when "0010100110000001" => data <= "111111";
				when "0010100110000100" => data <= "111111";
				when "0010100110000101" => data <= "010010";
				when "0010100110000110" => data <= "010010";
				when "0010100110000111" => data <= "010010";
				when "0010100110001000" => data <= "111111";
				when "0010101000011011" => data <= "111111";
				when "0010101000011100" => data <= "010010";
				when "0010101000011101" => data <= "010010";
				when "0010101000011110" => data <= "111111";
				when "0010101000100011" => data <= "111111";
				when "0010101000100100" => data <= "010010";
				when "0010101000100101" => data <= "010010";
				when "0010101000100110" => data <= "111111";
				when "0010101000101011" => data <= "111111";
				when "0010101000101100" => data <= "010010";
				when "0010101000101101" => data <= "010010";
				when "0010101000101110" => data <= "111111";
				when "0010101000110011" => data <= "111111";
				when "0010101000110100" => data <= "010010";
				when "0010101000110101" => data <= "010010";
				when "0010101000110110" => data <= "111111";
				when "0010101000111011" => data <= "111111";
				when "0010101000111100" => data <= "010010";
				when "0010101000111101" => data <= "010010";
				when "0010101000111110" => data <= "111111";
				when "0010101001000011" => data <= "111111";
				when "0010101001000100" => data <= "010010";
				when "0010101001000101" => data <= "010010";
				when "0010101001000110" => data <= "111111";
				when "0010101001001111" => data <= "111111";
				when "0010101001010000" => data <= "010010";
				when "0010101001010001" => data <= "010010";
				when "0010101001010010" => data <= "111111";
				when "0010101001011100" => data <= "111111";
				when "0010101001011101" => data <= "010010";
				when "0010101001011110" => data <= "010010";
				when "0010101001011111" => data <= "111111";
				when "0010101001100100" => data <= "111111";
				when "0010101001100101" => data <= "010010";
				when "0010101001100110" => data <= "010010";
				when "0010101001100111" => data <= "111111";
				when "0010101001101100" => data <= "111111";
				when "0010101001101101" => data <= "010010";
				when "0010101001101110" => data <= "010010";
				when "0010101001101111" => data <= "111111";
				when "0010101001110100" => data <= "111111";
				when "0010101001110101" => data <= "010010";
				when "0010101001110110" => data <= "010010";
				when "0010101001110111" => data <= "111111";
				when "0010101001111101" => data <= "111111";
				when "0010101001111110" => data <= "010010";
				when "0010101001111111" => data <= "010010";
				when "0010101010000000" => data <= "010010";
				when "0010101010000001" => data <= "010010";
				when "0010101010000010" => data <= "111111";
				when "0010101010000011" => data <= "111111";
				when "0010101010000100" => data <= "010010";
				when "0010101010000101" => data <= "010010";
				when "0010101010000110" => data <= "010010";
				when "0010101010000111" => data <= "010010";
				when "0010101010001000" => data <= "111111";
				when "0010101100011011" => data <= "111111";
				when "0010101100011100" => data <= "100010";
				when "0010101100011101" => data <= "100010";
				when "0010101100011110" => data <= "111111";
				when "0010101100100011" => data <= "111111";
				when "0010101100100100" => data <= "100010";
				when "0010101100100101" => data <= "100010";
				when "0010101100100110" => data <= "111111";
				when "0010101100101011" => data <= "111111";
				when "0010101100101100" => data <= "100010";
				when "0010101100101101" => data <= "100010";
				when "0010101100101110" => data <= "111111";
				when "0010101100110011" => data <= "111111";
				when "0010101100110100" => data <= "100010";
				when "0010101100110101" => data <= "100010";
				when "0010101100110110" => data <= "111111";
				when "0010101100111011" => data <= "111111";
				when "0010101100111100" => data <= "100010";
				when "0010101100111101" => data <= "100010";
				when "0010101100111110" => data <= "111111";
				when "0010101101000011" => data <= "111111";
				when "0010101101000100" => data <= "100010";
				when "0010101101000101" => data <= "100010";
				when "0010101101000110" => data <= "111111";
				when "0010101101001111" => data <= "111111";
				when "0010101101010000" => data <= "010010";
				when "0010101101010001" => data <= "010010";
				when "0010101101010010" => data <= "111111";
				when "0010101101011100" => data <= "111111";
				when "0010101101011101" => data <= "100010";
				when "0010101101011110" => data <= "100010";
				when "0010101101011111" => data <= "111111";
				when "0010101101100100" => data <= "111111";
				when "0010101101100101" => data <= "100010";
				when "0010101101100110" => data <= "100010";
				when "0010101101100111" => data <= "111111";
				when "0010101101101100" => data <= "111111";
				when "0010101101101101" => data <= "100010";
				when "0010101101101110" => data <= "100010";
				when "0010101101101111" => data <= "111111";
				when "0010101101110100" => data <= "111111";
				when "0010101101110101" => data <= "100010";
				when "0010101101110110" => data <= "100010";
				when "0010101101110111" => data <= "111111";
				when "0010101101111101" => data <= "111111";
				when "0010101101111110" => data <= "010010";
				when "0010101101111111" => data <= "010010";
				when "0010101110000000" => data <= "010010";
				when "0010101110000001" => data <= "010010";
				when "0010101110000010" => data <= "010010";
				when "0010101110000011" => data <= "010010";
				when "0010101110000100" => data <= "010010";
				when "0010101110000101" => data <= "010010";
				when "0010101110000110" => data <= "010010";
				when "0010101110000111" => data <= "010010";
				when "0010101110001000" => data <= "111111";
				when "0010110000011011" => data <= "111111";
				when "0010110000011100" => data <= "100010";
				when "0010110000011101" => data <= "100010";
				when "0010110000011110" => data <= "111111";
				when "0010110000100011" => data <= "111111";
				when "0010110000100100" => data <= "100010";
				when "0010110000100101" => data <= "100010";
				when "0010110000100110" => data <= "111111";
				when "0010110000101011" => data <= "111111";
				when "0010110000101100" => data <= "100010";
				when "0010110000101101" => data <= "100010";
				when "0010110000101110" => data <= "111111";
				when "0010110000110011" => data <= "111111";
				when "0010110000110100" => data <= "100010";
				when "0010110000110101" => data <= "100010";
				when "0010110000110110" => data <= "111111";
				when "0010110000111011" => data <= "111111";
				when "0010110000111100" => data <= "100010";
				when "0010110000111101" => data <= "100010";
				when "0010110000111110" => data <= "100010";
				when "0010110000111111" => data <= "111111";
				when "0010110001000010" => data <= "111111";
				when "0010110001000011" => data <= "100010";
				when "0010110001000100" => data <= "100010";
				when "0010110001000101" => data <= "100010";
				when "0010110001000110" => data <= "111111";
				when "0010110001001111" => data <= "111111";
				when "0010110001010000" => data <= "100010";
				when "0010110001010001" => data <= "100010";
				when "0010110001010010" => data <= "111111";
				when "0010110001011100" => data <= "111111";
				when "0010110001011101" => data <= "100010";
				when "0010110001011110" => data <= "100010";
				when "0010110001011111" => data <= "111111";
				when "0010110001100100" => data <= "111111";
				when "0010110001100101" => data <= "100010";
				when "0010110001100110" => data <= "100010";
				when "0010110001100111" => data <= "111111";
				when "0010110001101100" => data <= "111111";
				when "0010110001101101" => data <= "100010";
				when "0010110001101110" => data <= "100010";
				when "0010110001101111" => data <= "100010";
				when "0010110001110000" => data <= "111111";
				when "0010110001110011" => data <= "111111";
				when "0010110001110100" => data <= "111111";
				when "0010110001110101" => data <= "100010";
				when "0010110001110110" => data <= "100010";
				when "0010110001110111" => data <= "111111";
				when "0010110001111101" => data <= "111111";
				when "0010110001111110" => data <= "010010";
				when "0010110001111111" => data <= "010010";
				when "0010110010000000" => data <= "010010";
				when "0010110010000001" => data <= "111111";
				when "0010110010000010" => data <= "010010";
				when "0010110010000011" => data <= "010010";
				when "0010110010000100" => data <= "111111";
				when "0010110010000101" => data <= "010010";
				when "0010110010000110" => data <= "010010";
				when "0010110010000111" => data <= "010010";
				when "0010110010001000" => data <= "111111";
				when "0010110100011011" => data <= "111111";
				when "0010110100011100" => data <= "100010";
				when "0010110100011101" => data <= "100010";
				when "0010110100011110" => data <= "111111";
				when "0010110100100011" => data <= "111111";
				when "0010110100100100" => data <= "100010";
				when "0010110100100101" => data <= "100010";
				when "0010110100100110" => data <= "111111";
				when "0010110100101011" => data <= "111111";
				when "0010110100101100" => data <= "100010";
				when "0010110100101101" => data <= "100010";
				when "0010110100101110" => data <= "100010";
				when "0010110100101111" => data <= "111111";
				when "0010110100110000" => data <= "111111";
				when "0010110100110001" => data <= "111111";
				when "0010110100110010" => data <= "111111";
				when "0010110100110011" => data <= "100010";
				when "0010110100110100" => data <= "100010";
				when "0010110100110101" => data <= "100010";
				when "0010110100110110" => data <= "111111";
				when "0010110100111100" => data <= "111111";
				when "0010110100111101" => data <= "100010";
				when "0010110100111110" => data <= "100010";
				when "0010110100111111" => data <= "100010";
				when "0010110101000000" => data <= "111111";
				when "0010110101000001" => data <= "111111";
				when "0010110101000010" => data <= "100010";
				when "0010110101000011" => data <= "100010";
				when "0010110101000100" => data <= "100010";
				when "0010110101000101" => data <= "111111";
				when "0010110101001111" => data <= "111111";
				when "0010110101010000" => data <= "100010";
				when "0010110101010001" => data <= "100010";
				when "0010110101010010" => data <= "111111";
				when "0010110101011100" => data <= "111111";
				when "0010110101011101" => data <= "100010";
				when "0010110101011110" => data <= "100010";
				when "0010110101011111" => data <= "100010";
				when "0010110101100000" => data <= "111111";
				when "0010110101100001" => data <= "111111";
				when "0010110101100010" => data <= "111111";
				when "0010110101100011" => data <= "111111";
				when "0010110101100100" => data <= "100010";
				when "0010110101100101" => data <= "100010";
				when "0010110101100110" => data <= "100010";
				when "0010110101100111" => data <= "111111";
				when "0010110101101101" => data <= "111111";
				when "0010110101101110" => data <= "100010";
				when "0010110101101111" => data <= "100010";
				when "0010110101110000" => data <= "100010";
				when "0010110101110001" => data <= "111111";
				when "0010110101110010" => data <= "111111";
				when "0010110101110011" => data <= "100010";
				when "0010110101110100" => data <= "100010";
				when "0010110101110101" => data <= "100010";
				when "0010110101110110" => data <= "111111";
				when "0010110101111101" => data <= "111111";
				when "0010110101111110" => data <= "100010";
				when "0010110101111111" => data <= "100010";
				when "0010110110000000" => data <= "111111";
				when "0010110110000010" => data <= "111111";
				when "0010110110000011" => data <= "111111";
				when "0010110110000101" => data <= "111111";
				when "0010110110000110" => data <= "100010";
				when "0010110110000111" => data <= "100010";
				when "0010110110001000" => data <= "111111";
				when "0010111000011011" => data <= "111111";
				when "0010111000011100" => data <= "100010";
				when "0010111000011101" => data <= "100010";
				when "0010111000011110" => data <= "111111";
				when "0010111000011111" => data <= "111111";
				when "0010111000100000" => data <= "111111";
				when "0010111000100001" => data <= "111111";
				when "0010111000100010" => data <= "111111";
				when "0010111000100011" => data <= "111111";
				when "0010111000100100" => data <= "100010";
				when "0010111000100101" => data <= "100010";
				when "0010111000100110" => data <= "111111";
				when "0010111000101011" => data <= "111111";
				when "0010111000101100" => data <= "100010";
				when "0010111000101101" => data <= "100010";
				when "0010111000101110" => data <= "100010";
				when "0010111000101111" => data <= "100010";
				when "0010111000110000" => data <= "100010";
				when "0010111000110001" => data <= "100010";
				when "0010111000110010" => data <= "100010";
				when "0010111000110011" => data <= "100010";
				when "0010111000110100" => data <= "100010";
				when "0010111000110101" => data <= "100010";
				when "0010111000110110" => data <= "111111";
				when "0010111000111101" => data <= "111111";
				when "0010111000111110" => data <= "100010";
				when "0010111000111111" => data <= "100010";
				when "0010111001000000" => data <= "100010";
				when "0010111001000001" => data <= "100010";
				when "0010111001000010" => data <= "100010";
				when "0010111001000011" => data <= "100010";
				when "0010111001000100" => data <= "111111";
				when "0010111001001111" => data <= "111111";
				when "0010111001010000" => data <= "100010";
				when "0010111001010001" => data <= "100010";
				when "0010111001010010" => data <= "111111";
				when "0010111001011100" => data <= "111111";
				when "0010111001011101" => data <= "100010";
				when "0010111001011110" => data <= "100010";
				when "0010111001011111" => data <= "100010";
				when "0010111001100000" => data <= "100010";
				when "0010111001100001" => data <= "100010";
				when "0010111001100010" => data <= "100010";
				when "0010111001100011" => data <= "100010";
				when "0010111001100100" => data <= "100010";
				when "0010111001100101" => data <= "100010";
				when "0010111001100110" => data <= "100010";
				when "0010111001100111" => data <= "111111";
				when "0010111001101110" => data <= "111111";
				when "0010111001101111" => data <= "100010";
				when "0010111001110000" => data <= "100010";
				when "0010111001110001" => data <= "100010";
				when "0010111001110010" => data <= "100010";
				when "0010111001110011" => data <= "100010";
				when "0010111001110100" => data <= "100010";
				when "0010111001110101" => data <= "111111";
				when "0010111001111101" => data <= "111111";
				when "0010111001111110" => data <= "100010";
				when "0010111001111111" => data <= "100010";
				when "0010111010000000" => data <= "111111";
				when "0010111010000101" => data <= "111111";
				when "0010111010000110" => data <= "100010";
				when "0010111010000111" => data <= "100010";
				when "0010111010001000" => data <= "111111";
				when "0010111100011011" => data <= "111111";
				when "0010111100011100" => data <= "100010";
				when "0010111100011101" => data <= "100010";
				when "0010111100011110" => data <= "100010";
				when "0010111100011111" => data <= "100010";
				when "0010111100100000" => data <= "100010";
				when "0010111100100001" => data <= "100010";
				when "0010111100100010" => data <= "100010";
				when "0010111100100011" => data <= "100010";
				when "0010111100100100" => data <= "100010";
				when "0010111100100101" => data <= "111111";
				when "0010111100101011" => data <= "111111";
				when "0010111100101100" => data <= "100010";
				when "0010111100101101" => data <= "100010";
				when "0010111100101110" => data <= "100010";
				when "0010111100101111" => data <= "100010";
				when "0010111100110000" => data <= "100010";
				when "0010111100110001" => data <= "100010";
				when "0010111100110010" => data <= "100010";
				when "0010111100110011" => data <= "100010";
				when "0010111100110100" => data <= "100010";
				when "0010111100110101" => data <= "100010";
				when "0010111100110110" => data <= "111111";
				when "0010111100111110" => data <= "111111";
				when "0010111100111111" => data <= "100010";
				when "0010111101000000" => data <= "100010";
				when "0010111101000001" => data <= "100010";
				when "0010111101000010" => data <= "100010";
				when "0010111101000011" => data <= "111111";
				when "0010111101001111" => data <= "111111";
				when "0010111101010000" => data <= "100010";
				when "0010111101010001" => data <= "100010";
				when "0010111101010010" => data <= "111111";
				when "0010111101011100" => data <= "111111";
				when "0010111101011101" => data <= "100010";
				when "0010111101011110" => data <= "100010";
				when "0010111101011111" => data <= "100010";
				when "0010111101100000" => data <= "100010";
				when "0010111101100001" => data <= "100010";
				when "0010111101100010" => data <= "100010";
				when "0010111101100011" => data <= "100010";
				when "0010111101100100" => data <= "100010";
				when "0010111101100101" => data <= "100010";
				when "0010111101100110" => data <= "100010";
				when "0010111101100111" => data <= "111111";
				when "0010111101101111" => data <= "111111";
				when "0010111101110000" => data <= "100010";
				when "0010111101110001" => data <= "100010";
				when "0010111101110010" => data <= "100010";
				when "0010111101110011" => data <= "100010";
				when "0010111101110100" => data <= "111111";
				when "0010111101111101" => data <= "111111";
				when "0010111101111110" => data <= "100010";
				when "0010111101111111" => data <= "100010";
				when "0010111110000000" => data <= "111111";
				when "0010111110000101" => data <= "111111";
				when "0010111110000110" => data <= "100010";
				when "0010111110000111" => data <= "100010";
				when "0010111110001000" => data <= "111111";
				when "0011000000011011" => data <= "111111";
				when "0011000000011100" => data <= "100010";
				when "0011000000011101" => data <= "100010";
				when "0011000000011110" => data <= "100010";
				when "0011000000011111" => data <= "100010";
				when "0011000000100000" => data <= "100010";
				when "0011000000100001" => data <= "100010";
				when "0011000000100010" => data <= "100010";
				when "0011000000100011" => data <= "100010";
				when "0011000000100100" => data <= "111111";
				when "0011000000101011" => data <= "111111";
				when "0011000000101100" => data <= "100010";
				when "0011000000101101" => data <= "100010";
				when "0011000000101110" => data <= "100010";
				when "0011000000101111" => data <= "111111";
				when "0011000000110000" => data <= "111111";
				when "0011000000110001" => data <= "111111";
				when "0011000000110010" => data <= "111111";
				when "0011000000110011" => data <= "100010";
				when "0011000000110100" => data <= "100010";
				when "0011000000110101" => data <= "100010";
				when "0011000000110110" => data <= "111111";
				when "0011000000111111" => data <= "111111";
				when "0011000001000000" => data <= "100010";
				when "0011000001000001" => data <= "100010";
				when "0011000001000010" => data <= "111111";
				when "0011000001001111" => data <= "111111";
				when "0011000001010000" => data <= "100010";
				when "0011000001010001" => data <= "100010";
				when "0011000001010010" => data <= "111111";
				when "0011000001011100" => data <= "111111";
				when "0011000001011101" => data <= "100010";
				when "0011000001011110" => data <= "100010";
				when "0011000001011111" => data <= "100010";
				when "0011000001100000" => data <= "111111";
				when "0011000001100001" => data <= "111111";
				when "0011000001100010" => data <= "111111";
				when "0011000001100011" => data <= "111111";
				when "0011000001100100" => data <= "100010";
				when "0011000001100101" => data <= "100010";
				when "0011000001100110" => data <= "100010";
				when "0011000001100111" => data <= "111111";
				when "0011000001110000" => data <= "111111";
				when "0011000001110001" => data <= "100010";
				when "0011000001110010" => data <= "100010";
				when "0011000001110011" => data <= "111111";
				when "0011000001111101" => data <= "111111";
				when "0011000001111110" => data <= "100010";
				when "0011000001111111" => data <= "100010";
				when "0011000010000000" => data <= "111111";
				when "0011000010000101" => data <= "111111";
				when "0011000010000110" => data <= "100010";
				when "0011000010000111" => data <= "100010";
				when "0011000010001000" => data <= "111111";
				when "0011000100011011" => data <= "111111";
				when "0011000100011100" => data <= "100010";
				when "0011000100011101" => data <= "100010";
				when "0011000100011110" => data <= "100010";
				when "0011000100011111" => data <= "111111";
				when "0011000100100000" => data <= "111111";
				when "0011000100100001" => data <= "111111";
				when "0011000100100010" => data <= "111111";
				when "0011000100100011" => data <= "100010";
				when "0011000100100100" => data <= "100010";
				when "0011000100100101" => data <= "111111";
				when "0011000100101011" => data <= "111111";
				when "0011000100101100" => data <= "100010";
				when "0011000100101101" => data <= "100010";
				when "0011000100101110" => data <= "111111";
				when "0011000100110011" => data <= "111111";
				when "0011000100110100" => data <= "100010";
				when "0011000100110101" => data <= "100010";
				when "0011000100110110" => data <= "111111";
				when "0011000100111111" => data <= "111111";
				when "0011000101000000" => data <= "100010";
				when "0011000101000001" => data <= "100010";
				when "0011000101000010" => data <= "111111";
				when "0011000101001111" => data <= "111111";
				when "0011000101010000" => data <= "100010";
				when "0011000101010001" => data <= "100010";
				when "0011000101010010" => data <= "111111";
				when "0011000101011100" => data <= "111111";
				when "0011000101011101" => data <= "100010";
				when "0011000101011110" => data <= "100010";
				when "0011000101011111" => data <= "111111";
				when "0011000101100100" => data <= "111111";
				when "0011000101100101" => data <= "100010";
				when "0011000101100110" => data <= "100010";
				when "0011000101100111" => data <= "111111";
				when "0011000101110000" => data <= "111111";
				when "0011000101110001" => data <= "100010";
				when "0011000101110010" => data <= "100010";
				when "0011000101110011" => data <= "111111";
				when "0011000101111101" => data <= "111111";
				when "0011000101111110" => data <= "100010";
				when "0011000101111111" => data <= "100010";
				when "0011000110000000" => data <= "111111";
				when "0011000110000101" => data <= "111111";
				when "0011000110000110" => data <= "100010";
				when "0011000110000111" => data <= "100010";
				when "0011000110001000" => data <= "111111";
				when "0011001000011011" => data <= "111111";
				when "0011001000011100" => data <= "100010";
				when "0011001000011101" => data <= "100010";
				when "0011001000011110" => data <= "111111";
				when "0011001000100011" => data <= "111111";
				when "0011001000100100" => data <= "100010";
				when "0011001000100101" => data <= "100010";
				when "0011001000100110" => data <= "111111";
				when "0011001000101011" => data <= "111111";
				when "0011001000101100" => data <= "100010";
				when "0011001000101101" => data <= "100010";
				when "0011001000101110" => data <= "111111";
				when "0011001000110011" => data <= "111111";
				when "0011001000110100" => data <= "100010";
				when "0011001000110101" => data <= "100010";
				when "0011001000110110" => data <= "111111";
				when "0011001000111111" => data <= "111111";
				when "0011001001000000" => data <= "100010";
				when "0011001001000001" => data <= "100010";
				when "0011001001000010" => data <= "111111";
				when "0011001001001111" => data <= "111111";
				when "0011001001010000" => data <= "100010";
				when "0011001001010001" => data <= "100010";
				when "0011001001010010" => data <= "111111";
				when "0011001001011100" => data <= "111111";
				when "0011001001011101" => data <= "100010";
				when "0011001001011110" => data <= "100010";
				when "0011001001011111" => data <= "111111";
				when "0011001001100100" => data <= "111111";
				when "0011001001100101" => data <= "100010";
				when "0011001001100110" => data <= "100010";
				when "0011001001100111" => data <= "111111";
				when "0011001001110000" => data <= "111111";
				when "0011001001110001" => data <= "100010";
				when "0011001001110010" => data <= "100010";
				when "0011001001110011" => data <= "111111";
				when "0011001001111101" => data <= "111111";
				when "0011001001111110" => data <= "100010";
				when "0011001001111111" => data <= "100010";
				when "0011001010000000" => data <= "111111";
				when "0011001010000101" => data <= "111111";
				when "0011001010000110" => data <= "100010";
				when "0011001010000111" => data <= "100010";
				when "0011001010001000" => data <= "111111";
				when "0011001100011011" => data <= "111111";
				when "0011001100011100" => data <= "100010";
				when "0011001100011101" => data <= "100010";
				when "0011001100011110" => data <= "111111";
				when "0011001100100011" => data <= "111111";
				when "0011001100100100" => data <= "100010";
				when "0011001100100101" => data <= "100010";
				when "0011001100100110" => data <= "111111";
				when "0011001100101011" => data <= "111111";
				when "0011001100101100" => data <= "100010";
				when "0011001100101101" => data <= "100010";
				when "0011001100101110" => data <= "111111";
				when "0011001100110011" => data <= "111111";
				when "0011001100110100" => data <= "100010";
				when "0011001100110101" => data <= "100010";
				when "0011001100110110" => data <= "111111";
				when "0011001100111111" => data <= "111111";
				when "0011001101000000" => data <= "100010";
				when "0011001101000001" => data <= "100010";
				when "0011001101000010" => data <= "111111";
				when "0011001101001111" => data <= "111111";
				when "0011001101010000" => data <= "100010";
				when "0011001101010001" => data <= "100010";
				when "0011001101010010" => data <= "111111";
				when "0011001101011100" => data <= "111111";
				when "0011001101011101" => data <= "100010";
				when "0011001101011110" => data <= "100010";
				when "0011001101011111" => data <= "111111";
				when "0011001101100100" => data <= "111111";
				when "0011001101100101" => data <= "100010";
				when "0011001101100110" => data <= "100010";
				when "0011001101100111" => data <= "111111";
				when "0011001101110000" => data <= "111111";
				when "0011001101110001" => data <= "100010";
				when "0011001101110010" => data <= "100010";
				when "0011001101110011" => data <= "111111";
				when "0011001101111101" => data <= "111111";
				when "0011001101111110" => data <= "100010";
				when "0011001101111111" => data <= "100010";
				when "0011001110000000" => data <= "111111";
				when "0011001110000101" => data <= "111111";
				when "0011001110000110" => data <= "100010";
				when "0011001110000111" => data <= "100010";
				when "0011001110001000" => data <= "111111";
				when "0011010000011011" => data <= "111111";
				when "0011010000011100" => data <= "100010";
				when "0011010000011101" => data <= "100010";
				when "0011010000011110" => data <= "111111";
				when "0011010000100011" => data <= "111111";
				when "0011010000100100" => data <= "100010";
				when "0011010000100101" => data <= "100010";
				when "0011010000100110" => data <= "111111";
				when "0011010000101011" => data <= "111111";
				when "0011010000101100" => data <= "100010";
				when "0011010000101101" => data <= "100010";
				when "0011010000101110" => data <= "111111";
				when "0011010000110011" => data <= "111111";
				when "0011010000110100" => data <= "100010";
				when "0011010000110101" => data <= "100010";
				when "0011010000110110" => data <= "111111";
				when "0011010000111111" => data <= "111111";
				when "0011010001000000" => data <= "100010";
				when "0011010001000001" => data <= "100010";
				when "0011010001000010" => data <= "111111";
				when "0011010001001111" => data <= "111111";
				when "0011010001010000" => data <= "100010";
				when "0011010001010001" => data <= "100010";
				when "0011010001010010" => data <= "111111";
				when "0011010001011100" => data <= "111111";
				when "0011010001011101" => data <= "100010";
				when "0011010001011110" => data <= "100010";
				when "0011010001011111" => data <= "111111";
				when "0011010001100100" => data <= "111111";
				when "0011010001100101" => data <= "100010";
				when "0011010001100110" => data <= "100010";
				when "0011010001100111" => data <= "111111";
				when "0011010001110000" => data <= "111111";
				when "0011010001110001" => data <= "110010";
				when "0011010001110010" => data <= "110010";
				when "0011010001110011" => data <= "111111";
				when "0011010001111101" => data <= "111111";
				when "0011010001111110" => data <= "110010";
				when "0011010001111111" => data <= "110010";
				when "0011010010000000" => data <= "111111";
				when "0011010010000101" => data <= "111111";
				when "0011010010000110" => data <= "110010";
				when "0011010010000111" => data <= "110010";
				when "0011010010001000" => data <= "111111";
				when "0011010100011011" => data <= "111111";
				when "0011010100011100" => data <= "110010";
				when "0011010100011101" => data <= "110010";
				when "0011010100011110" => data <= "111111";
				when "0011010100100011" => data <= "111111";
				when "0011010100100100" => data <= "110010";
				when "0011010100100101" => data <= "110010";
				when "0011010100100110" => data <= "111111";
				when "0011010100101011" => data <= "111111";
				when "0011010100101100" => data <= "110010";
				when "0011010100101101" => data <= "110010";
				when "0011010100101110" => data <= "111111";
				when "0011010100110011" => data <= "111111";
				when "0011010100110100" => data <= "110010";
				when "0011010100110101" => data <= "110010";
				when "0011010100110110" => data <= "111111";
				when "0011010100111111" => data <= "111111";
				when "0011010101000000" => data <= "110010";
				when "0011010101000001" => data <= "110010";
				when "0011010101000010" => data <= "111111";
				when "0011010101001111" => data <= "111111";
				when "0011010101010000" => data <= "110010";
				when "0011010101010001" => data <= "110010";
				when "0011010101010010" => data <= "111111";
				when "0011010101011100" => data <= "111111";
				when "0011010101011101" => data <= "110010";
				when "0011010101011110" => data <= "110010";
				when "0011010101011111" => data <= "111111";
				when "0011010101100100" => data <= "111111";
				when "0011010101100101" => data <= "110010";
				when "0011010101100110" => data <= "110010";
				when "0011010101100111" => data <= "111111";
				when "0011010101110000" => data <= "111111";
				when "0011010101110001" => data <= "110010";
				when "0011010101110010" => data <= "110010";
				when "0011010101110011" => data <= "111111";
				when "0011010101111101" => data <= "111111";
				when "0011010101111110" => data <= "110010";
				when "0011010101111111" => data <= "110010";
				when "0011010110000000" => data <= "111111";
				when "0011010110000101" => data <= "111111";
				when "0011010110000110" => data <= "110010";
				when "0011010110000111" => data <= "110010";
				when "0011010110001000" => data <= "111111";
				when "0011011000011011" => data <= "111111";
				when "0011011000011100" => data <= "110010";
				when "0011011000011101" => data <= "110010";
				when "0011011000011110" => data <= "111111";
				when "0011011000100011" => data <= "111111";
				when "0011011000100100" => data <= "110010";
				when "0011011000100101" => data <= "110010";
				when "0011011000100110" => data <= "111111";
				when "0011011000101011" => data <= "111111";
				when "0011011000101100" => data <= "110010";
				when "0011011000101101" => data <= "110010";
				when "0011011000101110" => data <= "111111";
				when "0011011000110011" => data <= "111111";
				when "0011011000110100" => data <= "110010";
				when "0011011000110101" => data <= "110010";
				when "0011011000110110" => data <= "111111";
				when "0011011000111111" => data <= "111111";
				when "0011011001000000" => data <= "110010";
				when "0011011001000001" => data <= "110010";
				when "0011011001000010" => data <= "111111";
				when "0011011001001111" => data <= "111111";
				when "0011011001010000" => data <= "110010";
				when "0011011001010001" => data <= "110010";
				when "0011011001010010" => data <= "111111";
				when "0011011001011100" => data <= "111111";
				when "0011011001011101" => data <= "110010";
				when "0011011001011110" => data <= "110010";
				when "0011011001011111" => data <= "111111";
				when "0011011001100100" => data <= "111111";
				when "0011011001100101" => data <= "110010";
				when "0011011001100110" => data <= "110010";
				when "0011011001100111" => data <= "111111";
				when "0011011001110000" => data <= "111111";
				when "0011011001110001" => data <= "110010";
				when "0011011001110010" => data <= "110010";
				when "0011011001110011" => data <= "111111";
				when "0011011001111101" => data <= "111111";
				when "0011011001111110" => data <= "110010";
				when "0011011001111111" => data <= "110010";
				when "0011011010000000" => data <= "111111";
				when "0011011010000101" => data <= "111111";
				when "0011011010000110" => data <= "110010";
				when "0011011010000111" => data <= "110010";
				when "0011011010001000" => data <= "111111";
				when "0011011100011011" => data <= "111111";
				when "0011011100011100" => data <= "110010";
				when "0011011100011101" => data <= "110010";
				when "0011011100011110" => data <= "111111";
				when "0011011100100011" => data <= "111111";
				when "0011011100100100" => data <= "110010";
				when "0011011100100101" => data <= "110010";
				when "0011011100100110" => data <= "111111";
				when "0011011100101011" => data <= "111111";
				when "0011011100101100" => data <= "110010";
				when "0011011100101101" => data <= "110010";
				when "0011011100101110" => data <= "111111";
				when "0011011100110011" => data <= "111111";
				when "0011011100110100" => data <= "110010";
				when "0011011100110101" => data <= "110010";
				when "0011011100110110" => data <= "111111";
				when "0011011100111111" => data <= "111111";
				when "0011011101000000" => data <= "110010";
				when "0011011101000001" => data <= "110010";
				when "0011011101000010" => data <= "111111";
				when "0011011101001111" => data <= "111111";
				when "0011011101010000" => data <= "110010";
				when "0011011101010001" => data <= "110010";
				when "0011011101010010" => data <= "111111";
				when "0011011101011100" => data <= "111111";
				when "0011011101011101" => data <= "110010";
				when "0011011101011110" => data <= "110010";
				when "0011011101011111" => data <= "111111";
				when "0011011101100100" => data <= "111111";
				when "0011011101100101" => data <= "110010";
				when "0011011101100110" => data <= "110010";
				when "0011011101100111" => data <= "111111";
				when "0011011101110000" => data <= "111111";
				when "0011011101110001" => data <= "110010";
				when "0011011101110010" => data <= "110010";
				when "0011011101110011" => data <= "111111";
				when "0011011101111101" => data <= "111111";
				when "0011011101111110" => data <= "110010";
				when "0011011101111111" => data <= "110010";
				when "0011011110000000" => data <= "111111";
				when "0011011110000101" => data <= "111111";
				when "0011011110000110" => data <= "110010";
				when "0011011110000111" => data <= "110010";
				when "0011011110001000" => data <= "111111";
				when "0011100000011100" => data <= "111111";
				when "0011100000011101" => data <= "111111";
				when "0011100000100100" => data <= "111111";
				when "0011100000100101" => data <= "111111";
				when "0011100000101100" => data <= "111111";
				when "0011100000101101" => data <= "111111";
				when "0011100000110100" => data <= "111111";
				when "0011100000110101" => data <= "111111";
				when "0011100001000000" => data <= "111111";
				when "0011100001000001" => data <= "111111";
				when "0011100001010000" => data <= "111111";
				when "0011100001010001" => data <= "111111";
				when "0011100001011101" => data <= "111111";
				when "0011100001011110" => data <= "111111";
				when "0011100001100101" => data <= "111111";
				when "0011100001100110" => data <= "111111";
				when "0011100001110001" => data <= "111111";
				when "0011100001110010" => data <= "111111";
				when "0011100001111110" => data <= "111111";
				when "0011100001111111" => data <= "111111";
				when "0011100010000110" => data <= "111111";
				when "0011100010000111" => data <= "111111";
				when "0011101101000000" => data <= "100010";
				when "0011101101000001" => data <= "100010";
				when "0011101101000010" => data <= "100010";
				when "0011101101000011" => data <= "100010";
				when "0011101101000100" => data <= "100010";
				when "0011101101100010" => data <= "100010";
				when "0011110001000000" => data <= "100010";
				when "0011110001000001" => data <= "100010";
				when "0011110001000010" => data <= "100010";
				when "0011110001000011" => data <= "100010";
				when "0011110001000100" => data <= "100010";
				when "0011110001100010" => data <= "100010";
				when "0011110101000000" => data <= "100010";
				when "0011110101000100" => data <= "100010";
				when "0011110101000101" => data <= "100010";
				when "0011110101100010" => data <= "100010";
				when "0011111001000000" => data <= "100010";
				when "0011111001000100" => data <= "100010";
				when "0011111001000101" => data <= "100010";
				when "0011111001001101" => data <= "100010";
				when "0011111001001110" => data <= "100010";
				when "0011111001001111" => data <= "100010";
				when "0011111001010000" => data <= "100010";
				when "0011111001010001" => data <= "100010";
				when "0011111001010010" => data <= "100010";
				when "0011111001010011" => data <= "100010";
				when "0011111001010100" => data <= "100010";
				when "0011111001010101" => data <= "100010";
				when "0011111001010110" => data <= "100010";
				when "0011111001100010" => data <= "100010";
				when "0011111101000000" => data <= "100010";
				when "0011111101000101" => data <= "100010";
				when "0011111101000110" => data <= "100010";
				when "0011111101001101" => data <= "100010";
				when "0011111101010110" => data <= "100010";
				when "0011111101100010" => data <= "100010";
				when "0100000001000000" => data <= "100010";
				when "0100000001000101" => data <= "100010";
				when "0100000001000110" => data <= "100010";
				when "0100000001001101" => data <= "100010";
				when "0100000001001110" => data <= "100010";
				when "0100000001001111" => data <= "100010";
				when "0100000001010000" => data <= "100010";
				when "0100000001010001" => data <= "100010";
				when "0100000001010010" => data <= "100010";
				when "0100000001010011" => data <= "100010";
				when "0100000001010100" => data <= "100010";
				when "0100000001010101" => data <= "100010";
				when "0100000001010110" => data <= "100010";
				when "0100000001100010" => data <= "100010";
				when "0100000101000000" => data <= "100010";
				when "0100000101000101" => data <= "100010";
				when "0100000101001101" => data <= "100010";
				when "0100000101010110" => data <= "100010";
				when "0100000101100010" => data <= "100010";
				when "0100001001000000" => data <= "100010";
				when "0100001001000100" => data <= "010010";
				when "0100001001001101" => data <= "100010";
				when "0100001001010110" => data <= "100010";
				when "0100001001100010" => data <= "100010";
				when "0100001101000000" => data <= "100010";
				when "0100001101001101" => data <= "100010";
				when "0100001101010110" => data <= "100010";
				when "0100001101100010" => data <= "100010";
				when "0100010001000000" => data <= "100010";
				when "0100010001001101" => data <= "100010";
				when "0100010001010110" => data <= "100010";
				when "0100010001011101" => data <= "100010";
				when "0100010001011110" => data <= "100010";
				when "0100010001011111" => data <= "100010";
				when "0100010001100000" => data <= "100010";
				when "0100010001100001" => data <= "100010";
				when "0100010001100010" => data <= "100010";
				when "0100010100111100" => data <= "100010";
				when "0100010100111101" => data <= "100010";
				when "0100010100111110" => data <= "100010";
				when "0100010100111111" => data <= "100010";
				when "0100010101000000" => data <= "100010";
				when "0100010101001101" => data <= "100010";
				when "0100010101010110" => data <= "100010";
				when "0100010101011100" => data <= "100010";
				when "0100010101011101" => data <= "100010";
				when "0100010101011110" => data <= "100010";
				when "0100010101011111" => data <= "100010";
				when "0100010101100000" => data <= "100010";
				when "0100010101100001" => data <= "100010";
				when "0100010101100010" => data <= "100010";
				when "0100011000111011" => data <= "100010";
				when "0100011000111100" => data <= "100010";
				when "0100011000111101" => data <= "100010";
				when "0100011000111110" => data <= "100010";
				when "0100011000111111" => data <= "100010";
				when "0100011001000000" => data <= "100010";
				when "0100011001001001" => data <= "100010";
				when "0100011001001010" => data <= "100010";
				when "0100011001001011" => data <= "100010";
				when "0100011001001100" => data <= "100010";
				when "0100011001001101" => data <= "100010";
				when "0100011001010010" => data <= "100010";
				when "0100011001010011" => data <= "100010";
				when "0100011001010100" => data <= "100010";
				when "0100011001010101" => data <= "100010";
				when "0100011001010110" => data <= "100010";
				when "0100011001011100" => data <= "100010";
				when "0100011001011101" => data <= "111111";
				when "0100011001011110" => data <= "100010";
				when "0100011001011111" => data <= "100010";
				when "0100011001100000" => data <= "100010";
				when "0100011001100001" => data <= "100010";
				when "0100011001100010" => data <= "100010";
				when "0100011100111011" => data <= "100010";
				when "0100011100111100" => data <= "111111";
				when "0100011100111101" => data <= "100010";
				when "0100011100111110" => data <= "100010";
				when "0100011100111111" => data <= "100010";
				when "0100011101000000" => data <= "100010";
				when "0100011101001000" => data <= "100010";
				when "0100011101001001" => data <= "100010";
				when "0100011101001010" => data <= "100010";
				when "0100011101001011" => data <= "100010";
				when "0100011101001100" => data <= "100010";
				when "0100011101001101" => data <= "100010";
				when "0100011101010001" => data <= "100010";
				when "0100011101010010" => data <= "100010";
				when "0100011101010011" => data <= "100010";
				when "0100011101010100" => data <= "100010";
				when "0100011101010101" => data <= "100010";
				when "0100011101010110" => data <= "100010";
				when "0100011101011100" => data <= "100010";
				when "0100011101011101" => data <= "100010";
				when "0100011101011110" => data <= "100010";
				when "0100011101011111" => data <= "100010";
				when "0100011101100000" => data <= "100010";
				when "0100011101100001" => data <= "100010";
				when "0100011101100010" => data <= "100010";
				when "0100100000111011" => data <= "110010";
				when "0100100000111100" => data <= "110010";
				when "0100100000111101" => data <= "100010";
				when "0100100000111110" => data <= "100010";
				when "0100100000111111" => data <= "110010";
				when "0100100001000000" => data <= "110010";
				when "0100100001001000" => data <= "100010";
				when "0100100001001001" => data <= "111111";
				when "0100100001001010" => data <= "100010";
				when "0100100001001011" => data <= "100010";
				when "0100100001001100" => data <= "100010";
				when "0100100001001101" => data <= "100010";
				when "0100100001010001" => data <= "100010";
				when "0100100001010010" => data <= "111111";
				when "0100100001010011" => data <= "100010";
				when "0100100001010100" => data <= "100010";
				when "0100100001010101" => data <= "100010";
				when "0100100001010110" => data <= "100010";
				when "0100100001011100" => data <= "110010";
				when "0100100001011101" => data <= "110010";
				when "0100100001011110" => data <= "100010";
				when "0100100001011111" => data <= "100010";
				when "0100100001100000" => data <= "100010";
				when "0100100001100001" => data <= "110010";
				when "0100100001100010" => data <= "110010";
				when "0100100100111011" => data <= "100010";
				when "0100100100111100" => data <= "110010";
				when "0100100100111101" => data <= "110010";
				when "0100100100111110" => data <= "110010";
				when "0100100100111111" => data <= "110010";
				when "0100100101000000" => data <= "100010";
				when "0100100101001000" => data <= "110010";
				when "0100100101001001" => data <= "110010";
				when "0100100101001010" => data <= "100010";
				when "0100100101001011" => data <= "100010";
				when "0100100101001100" => data <= "110010";
				when "0100100101001101" => data <= "110010";
				when "0100100101010001" => data <= "110010";
				when "0100100101010010" => data <= "110010";
				when "0100100101010011" => data <= "100010";
				when "0100100101010100" => data <= "100010";
				when "0100100101010101" => data <= "110010";
				when "0100100101010110" => data <= "110010";
				when "0100100101011100" => data <= "100010";
				when "0100100101011101" => data <= "110010";
				when "0100100101011110" => data <= "110010";
				when "0100100101011111" => data <= "100010";
				when "0100100101100000" => data <= "110010";
				when "0100100101100001" => data <= "110010";
				when "0100100101100010" => data <= "100010";
				when "0100101000111011" => data <= "100010";
				when "0100101000111100" => data <= "100010";
				when "0100101000111101" => data <= "110010";
				when "0100101000111110" => data <= "110010";
				when "0100101000111111" => data <= "100010";
				when "0100101001000000" => data <= "100010";
				when "0100101001001000" => data <= "100010";
				when "0100101001001001" => data <= "110010";
				when "0100101001001010" => data <= "110010";
				when "0100101001001011" => data <= "110010";
				when "0100101001001100" => data <= "110010";
				when "0100101001001101" => data <= "100010";
				when "0100101001010001" => data <= "100010";
				when "0100101001010010" => data <= "110010";
				when "0100101001010011" => data <= "110010";
				when "0100101001010100" => data <= "110010";
				when "0100101001010101" => data <= "110010";
				when "0100101001010110" => data <= "100010";
				when "0100101001011100" => data <= "100010";
				when "0100101001011101" => data <= "100010";
				when "0100101001011110" => data <= "110010";
				when "0100101001011111" => data <= "110010";
				when "0100101001100000" => data <= "110010";
				when "0100101001100001" => data <= "100010";
				when "0100101001100010" => data <= "100010";
				when "0100101100111100" => data <= "100010";
				when "0100101100111101" => data <= "100010";
				when "0100101100111110" => data <= "100010";
				when "0100101100111111" => data <= "100010";
				when "0100101101001000" => data <= "100010";
				when "0100101101001001" => data <= "100010";
				when "0100101101001010" => data <= "110010";
				when "0100101101001011" => data <= "110010";
				when "0100101101001100" => data <= "100010";
				when "0100101101001101" => data <= "100010";
				when "0100101101010001" => data <= "100010";
				when "0100101101010010" => data <= "100010";
				when "0100101101010011" => data <= "110010";
				when "0100101101010100" => data <= "110010";
				when "0100101101010101" => data <= "100010";
				when "0100101101010110" => data <= "100010";
				when "0100101101011101" => data <= "100010";
				when "0100101101011110" => data <= "100010";
				when "0100101101011111" => data <= "100010";
				when "0100101101100000" => data <= "100010";
				when "0100101101100001" => data <= "100010";
				when "0100110001001001" => data <= "100010";
				when "0100110001001010" => data <= "100010";
				when "0100110001001011" => data <= "100010";
				when "0100110001001100" => data <= "100010";
				when "0100110001010010" => data <= "100010";
				when "0100110001010011" => data <= "100010";
				when "0100110001010100" => data <= "100010";
				when "0100110001010101" => data <= "100010";
				when "0101010100011111" => data <= "111111";
				when "0101010100100000" => data <= "111111";
				when "0101010100100001" => data <= "111111";
				when "0101010100100010" => data <= "111111";
				when "0101010100100011" => data <= "111111";
				when "0101010100101000" => data <= "111111";
				when "0101010100101001" => data <= "111111";
				when "0101010100101010" => data <= "111111";
				when "0101010100101011" => data <= "111111";
				when "0101010100101100" => data <= "111111";
				when "0101010100101101" => data <= "111111";
				when "0101010100110001" => data <= "111111";
				when "0101010100110010" => data <= "111111";
				when "0101010100110011" => data <= "111111";
				when "0101010100110100" => data <= "111111";
				when "0101010100110101" => data <= "111111";
				when "0101010100110110" => data <= "111111";
				when "0101010100110111" => data <= "111111";
				when "0101010100111011" => data <= "111111";
				when "0101010100111100" => data <= "111111";
				when "0101010100111101" => data <= "111111";
				when "0101010100111110" => data <= "111111";
				when "0101010100111111" => data <= "111111";
				when "0101010101000000" => data <= "111111";
				when "0101010101000101" => data <= "111111";
				when "0101010101000110" => data <= "111111";
				when "0101010101000111" => data <= "111111";
				when "0101010101001000" => data <= "111111";
				when "0101010101001001" => data <= "111111";
				when "0101010101001010" => data <= "111111";
				when "0101010101001011" => data <= "111111";
				when "0101010101010110" => data <= "111111";
				when "0101010101010111" => data <= "111111";
				when "0101010101011000" => data <= "111111";
				when "0101010101011001" => data <= "111111";
				when "0101010101011010" => data <= "111111";
				when "0101010101011011" => data <= "111111";
				when "0101010101011100" => data <= "111111";
				when "0101010101011111" => data <= "111111";
				when "0101010101100000" => data <= "111111";
				when "0101010101100001" => data <= "111111";
				when "0101010101100010" => data <= "111111";
				when "0101010101100011" => data <= "111111";
				when "0101010101100100" => data <= "111111";
				when "0101010101100101" => data <= "111111";
				when "0101010101100110" => data <= "111111";
				when "0101010101101011" => data <= "111111";
				when "0101010101101100" => data <= "111111";
				when "0101010101110101" => data <= "111111";
				when "0101010101110110" => data <= "111111";
				when "0101010101110111" => data <= "111111";
				when "0101010101111000" => data <= "111111";
				when "0101010101111001" => data <= "111111";
				when "0101010101111010" => data <= "111111";
				when "0101010101111110" => data <= "111111";
				when "0101010101111111" => data <= "111111";
				when "0101010110000000" => data <= "111111";
				when "0101010110000001" => data <= "111111";
				when "0101010110000010" => data <= "111111";
				when "0101010110000011" => data <= "111111";
				when "0101010110000100" => data <= "111111";
				when "0101010110000101" => data <= "111111";
				when "0101011000011110" => data <= "111111";
				when "0101011000011111" => data <= "111111";
				when "0101011000100000" => data <= "111111";
				when "0101011000100001" => data <= "111111";
				when "0101011000100010" => data <= "111111";
				when "0101011000100011" => data <= "111111";
				when "0101011000100111" => data <= "111111";
				when "0101011000101000" => data <= "111111";
				when "0101011000101001" => data <= "111111";
				when "0101011000101010" => data <= "111111";
				when "0101011000101011" => data <= "111111";
				when "0101011000101100" => data <= "111111";
				when "0101011000101101" => data <= "111111";
				when "0101011000101110" => data <= "111111";
				when "0101011000110001" => data <= "111111";
				when "0101011000110010" => data <= "111111";
				when "0101011000110011" => data <= "111111";
				when "0101011000110100" => data <= "111111";
				when "0101011000110101" => data <= "111111";
				when "0101011000110110" => data <= "111111";
				when "0101011000110111" => data <= "111111";
				when "0101011000111011" => data <= "111111";
				when "0101011000111100" => data <= "111111";
				when "0101011000111101" => data <= "111111";
				when "0101011000111110" => data <= "111111";
				when "0101011000111111" => data <= "111111";
				when "0101011001000000" => data <= "111111";
				when "0101011001000101" => data <= "111111";
				when "0101011001000110" => data <= "111111";
				when "0101011001000111" => data <= "111111";
				when "0101011001001000" => data <= "111111";
				when "0101011001001001" => data <= "111111";
				when "0101011001001010" => data <= "111111";
				when "0101011001001011" => data <= "111111";
				when "0101011001010110" => data <= "111111";
				when "0101011001010111" => data <= "111111";
				when "0101011001011000" => data <= "111111";
				when "0101011001011001" => data <= "111111";
				when "0101011001011010" => data <= "111111";
				when "0101011001011011" => data <= "111111";
				when "0101011001011100" => data <= "111111";
				when "0101011001011111" => data <= "111111";
				when "0101011001100000" => data <= "111111";
				when "0101011001100001" => data <= "111111";
				when "0101011001100010" => data <= "111111";
				when "0101011001100011" => data <= "111111";
				when "0101011001100100" => data <= "111111";
				when "0101011001100101" => data <= "111111";
				when "0101011001100110" => data <= "111111";
				when "0101011001101011" => data <= "111111";
				when "0101011001101100" => data <= "111111";
				when "0101011001110100" => data <= "111111";
				when "0101011001110101" => data <= "111111";
				when "0101011001110110" => data <= "111111";
				when "0101011001110111" => data <= "111111";
				when "0101011001111000" => data <= "111111";
				when "0101011001111001" => data <= "111111";
				when "0101011001111010" => data <= "111111";
				when "0101011001111011" => data <= "111111";
				when "0101011001111110" => data <= "111111";
				when "0101011001111111" => data <= "111111";
				when "0101011010000000" => data <= "111111";
				when "0101011010000001" => data <= "111111";
				when "0101011010000010" => data <= "111111";
				when "0101011010000011" => data <= "111111";
				when "0101011010000100" => data <= "111111";
				when "0101011010000101" => data <= "111111";
				when "0101011100011110" => data <= "111111";
				when "0101011100011111" => data <= "111111";
				when "0101011100100100" => data <= "111111";
				when "0101011100100101" => data <= "111111";
				when "0101011100100111" => data <= "111111";
				when "0101011100101000" => data <= "111111";
				when "0101011100101101" => data <= "111111";
				when "0101011100101110" => data <= "111111";
				when "0101011100110001" => data <= "111111";
				when "0101011100110010" => data <= "111111";
				when "0101011100111001" => data <= "111111";
				when "0101011100111010" => data <= "111111";
				when "0101011101000011" => data <= "111111";
				when "0101011101000100" => data <= "111111";
				when "0101011101010101" => data <= "111111";
				when "0101011101010110" => data <= "111111";
				when "0101011101100010" => data <= "111111";
				when "0101011101100011" => data <= "111111";
				when "0101011101101001" => data <= "111111";
				when "0101011101101010" => data <= "111111";
				when "0101011101101101" => data <= "111111";
				when "0101011101101110" => data <= "111111";
				when "0101011101110100" => data <= "111111";
				when "0101011101110101" => data <= "111111";
				when "0101011101111010" => data <= "111111";
				when "0101011101111011" => data <= "111111";
				when "0101011110000001" => data <= "111111";
				when "0101011110000010" => data <= "111111";
				when "0101100000011110" => data <= "111111";
				when "0101100000011111" => data <= "111111";
				when "0101100000100100" => data <= "111111";
				when "0101100000100101" => data <= "111111";
				when "0101100000100111" => data <= "111111";
				when "0101100000101000" => data <= "111111";
				when "0101100000101101" => data <= "111111";
				when "0101100000101110" => data <= "111111";
				when "0101100000110001" => data <= "111111";
				when "0101100000110010" => data <= "111111";
				when "0101100000111001" => data <= "111111";
				when "0101100000111010" => data <= "111111";
				when "0101100001000011" => data <= "111111";
				when "0101100001000100" => data <= "111111";
				when "0101100001010101" => data <= "111111";
				when "0101100001010110" => data <= "111111";
				when "0101100001100010" => data <= "111111";
				when "0101100001100011" => data <= "111111";
				when "0101100001101001" => data <= "111111";
				when "0101100001101010" => data <= "111111";
				when "0101100001101101" => data <= "111111";
				when "0101100001101110" => data <= "111111";
				when "0101100001110100" => data <= "111111";
				when "0101100001110101" => data <= "111111";
				when "0101100001111010" => data <= "111111";
				when "0101100001111011" => data <= "111111";
				when "0101100010000001" => data <= "111111";
				when "0101100010000010" => data <= "111111";
				when "0101100100011110" => data <= "111111";
				when "0101100100011111" => data <= "111111";
				when "0101100100100100" => data <= "111111";
				when "0101100100100101" => data <= "111111";
				when "0101100100100111" => data <= "111111";
				when "0101100100101000" => data <= "111111";
				when "0101100100101101" => data <= "111111";
				when "0101100100101110" => data <= "111111";
				when "0101100100110001" => data <= "111111";
				when "0101100100110010" => data <= "111111";
				when "0101100100111001" => data <= "111111";
				when "0101100100111010" => data <= "111111";
				when "0101100101000011" => data <= "111111";
				when "0101100101000100" => data <= "111111";
				when "0101100101010101" => data <= "111111";
				when "0101100101010110" => data <= "111111";
				when "0101100101100010" => data <= "111111";
				when "0101100101100011" => data <= "111111";
				when "0101100101100111" => data <= "111111";
				when "0101100101101000" => data <= "111111";
				when "0101100101101111" => data <= "111111";
				when "0101100101110000" => data <= "111111";
				when "0101100101110100" => data <= "111111";
				when "0101100101110101" => data <= "111111";
				when "0101100101111010" => data <= "111111";
				when "0101100101111011" => data <= "111111";
				when "0101100110000001" => data <= "111111";
				when "0101100110000010" => data <= "111111";
				when "0101101000011110" => data <= "111111";
				when "0101101000011111" => data <= "111111";
				when "0101101000100100" => data <= "111111";
				when "0101101000100101" => data <= "111111";
				when "0101101000100111" => data <= "111111";
				when "0101101000101000" => data <= "111111";
				when "0101101000101101" => data <= "111111";
				when "0101101000101110" => data <= "111111";
				when "0101101000110001" => data <= "111111";
				when "0101101000110010" => data <= "111111";
				when "0101101000111001" => data <= "111111";
				when "0101101000111010" => data <= "111111";
				when "0101101001000011" => data <= "111111";
				when "0101101001000100" => data <= "111111";
				when "0101101001010101" => data <= "111111";
				when "0101101001010110" => data <= "111111";
				when "0101101001100010" => data <= "111111";
				when "0101101001100011" => data <= "111111";
				when "0101101001100111" => data <= "111111";
				when "0101101001101000" => data <= "111111";
				when "0101101001101111" => data <= "111111";
				when "0101101001110000" => data <= "111111";
				when "0101101001110100" => data <= "111111";
				when "0101101001110101" => data <= "111111";
				when "0101101001111010" => data <= "111111";
				when "0101101001111011" => data <= "111111";
				when "0101101010000001" => data <= "111111";
				when "0101101010000010" => data <= "111111";
				when "0101101100011110" => data <= "111111";
				when "0101101100011111" => data <= "111111";
				when "0101101100100000" => data <= "111111";
				when "0101101100100001" => data <= "111111";
				when "0101101100100010" => data <= "111111";
				when "0101101100100011" => data <= "111111";
				when "0101101100100111" => data <= "111111";
				when "0101101100101000" => data <= "111111";
				when "0101101100101001" => data <= "111111";
				when "0101101100101010" => data <= "111111";
				when "0101101100101011" => data <= "111111";
				when "0101101100101100" => data <= "111111";
				when "0101101100110001" => data <= "111111";
				when "0101101100110010" => data <= "111111";
				when "0101101100110011" => data <= "111111";
				when "0101101100110100" => data <= "111111";
				when "0101101100110101" => data <= "111111";
				when "0101101100111001" => data <= "111111";
				when "0101101100111010" => data <= "111111";
				when "0101101100111011" => data <= "111111";
				when "0101101100111100" => data <= "111111";
				when "0101101100111101" => data <= "111111";
				when "0101101100111110" => data <= "111111";
				when "0101101100111111" => data <= "111111";
				when "0101101101000000" => data <= "111111";
				when "0101101101000011" => data <= "111111";
				when "0101101101000100" => data <= "111111";
				when "0101101101000101" => data <= "111111";
				when "0101101101000110" => data <= "111111";
				when "0101101101000111" => data <= "111111";
				when "0101101101001000" => data <= "111111";
				when "0101101101001001" => data <= "111111";
				when "0101101101001010" => data <= "111111";
				when "0101101101001011" => data <= "111111";
				when "0101101101010101" => data <= "111111";
				when "0101101101010110" => data <= "111111";
				when "0101101101010111" => data <= "111111";
				when "0101101101011000" => data <= "111111";
				when "0101101101011001" => data <= "111111";
				when "0101101101011010" => data <= "111111";
				when "0101101101011011" => data <= "111111";
				when "0101101101011100" => data <= "111111";
				when "0101101101100010" => data <= "111111";
				when "0101101101100011" => data <= "111111";
				when "0101101101100111" => data <= "111111";
				when "0101101101101000" => data <= "111111";
				when "0101101101101001" => data <= "111111";
				when "0101101101101010" => data <= "111111";
				when "0101101101101011" => data <= "111111";
				when "0101101101101100" => data <= "111111";
				when "0101101101101101" => data <= "111111";
				when "0101101101101110" => data <= "111111";
				when "0101101101101111" => data <= "111111";
				when "0101101101110000" => data <= "111111";
				when "0101101101110100" => data <= "111111";
				when "0101101101110101" => data <= "111111";
				when "0101101101110110" => data <= "111111";
				when "0101101101110111" => data <= "111111";
				when "0101101101111000" => data <= "111111";
				when "0101101101111001" => data <= "111111";
				when "0101101110000001" => data <= "111111";
				when "0101101110000010" => data <= "111111";
				when "0101110000011110" => data <= "111111";
				when "0101110000011111" => data <= "111111";
				when "0101110000100000" => data <= "111111";
				when "0101110000100001" => data <= "111111";
				when "0101110000100010" => data <= "111111";
				when "0101110000100011" => data <= "111111";
				when "0101110000100111" => data <= "111111";
				when "0101110000101000" => data <= "111111";
				when "0101110000101001" => data <= "111111";
				when "0101110000101010" => data <= "111111";
				when "0101110000101011" => data <= "111111";
				when "0101110000101100" => data <= "111111";
				when "0101110000101101" => data <= "111111";
				when "0101110000101110" => data <= "111111";
				when "0101110000110001" => data <= "111111";
				when "0101110000110010" => data <= "111111";
				when "0101110000110011" => data <= "111111";
				when "0101110000110100" => data <= "111111";
				when "0101110000110101" => data <= "111111";
				when "0101110000111011" => data <= "111111";
				when "0101110000111100" => data <= "111111";
				when "0101110000111101" => data <= "111111";
				when "0101110000111110" => data <= "111111";
				when "0101110000111111" => data <= "111111";
				when "0101110001000000" => data <= "111111";
				when "0101110001000001" => data <= "111111";
				when "0101110001000101" => data <= "111111";
				when "0101110001000110" => data <= "111111";
				when "0101110001000111" => data <= "111111";
				when "0101110001001000" => data <= "111111";
				when "0101110001001001" => data <= "111111";
				when "0101110001001010" => data <= "111111";
				when "0101110001001011" => data <= "111111";
				when "0101110001001100" => data <= "111111";
				when "0101110001010111" => data <= "111111";
				when "0101110001011000" => data <= "111111";
				when "0101110001011001" => data <= "111111";
				when "0101110001011010" => data <= "111111";
				when "0101110001011011" => data <= "111111";
				when "0101110001011100" => data <= "111111";
				when "0101110001011101" => data <= "111111";
				when "0101110001100010" => data <= "111111";
				when "0101110001100011" => data <= "111111";
				when "0101110001100111" => data <= "111111";
				when "0101110001101000" => data <= "111111";
				when "0101110001101001" => data <= "111111";
				when "0101110001101010" => data <= "111111";
				when "0101110001101011" => data <= "111111";
				when "0101110001101100" => data <= "111111";
				when "0101110001101101" => data <= "111111";
				when "0101110001101110" => data <= "111111";
				when "0101110001101111" => data <= "111111";
				when "0101110001110000" => data <= "111111";
				when "0101110001110100" => data <= "111111";
				when "0101110001110101" => data <= "111111";
				when "0101110001110110" => data <= "111111";
				when "0101110001110111" => data <= "111111";
				when "0101110001111000" => data <= "111111";
				when "0101110001111001" => data <= "111111";
				when "0101110001111010" => data <= "111111";
				when "0101110001111011" => data <= "111111";
				when "0101110010000001" => data <= "111111";
				when "0101110010000010" => data <= "111111";
				when "0101110100011110" => data <= "111111";
				when "0101110100011111" => data <= "111111";
				when "0101110100100111" => data <= "111111";
				when "0101110100101000" => data <= "111111";
				when "0101110100101101" => data <= "111111";
				when "0101110100101110" => data <= "111111";
				when "0101110100110001" => data <= "111111";
				when "0101110100110010" => data <= "111111";
				when "0101110101000000" => data <= "111111";
				when "0101110101000001" => data <= "111111";
				when "0101110101001011" => data <= "111111";
				when "0101110101001100" => data <= "111111";
				when "0101110101011100" => data <= "111111";
				when "0101110101011101" => data <= "111111";
				when "0101110101100010" => data <= "111111";
				when "0101110101100011" => data <= "111111";
				when "0101110101100111" => data <= "111111";
				when "0101110101101000" => data <= "111111";
				when "0101110101101111" => data <= "111111";
				when "0101110101110000" => data <= "111111";
				when "0101110101110100" => data <= "111111";
				when "0101110101110101" => data <= "111111";
				when "0101110101111010" => data <= "111111";
				when "0101110101111011" => data <= "111111";
				when "0101110110000001" => data <= "111111";
				when "0101110110000010" => data <= "111111";
				when "0101111000011110" => data <= "111111";
				when "0101111000011111" => data <= "111111";
				when "0101111000100111" => data <= "111111";
				when "0101111000101000" => data <= "111111";
				when "0101111000101101" => data <= "111111";
				when "0101111000101110" => data <= "111111";
				when "0101111000110001" => data <= "111111";
				when "0101111000110010" => data <= "111111";
				when "0101111001000000" => data <= "111111";
				when "0101111001000001" => data <= "111111";
				when "0101111001001011" => data <= "111111";
				when "0101111001001100" => data <= "111111";
				when "0101111001011100" => data <= "111111";
				when "0101111001011101" => data <= "111111";
				when "0101111001100010" => data <= "111111";
				when "0101111001100011" => data <= "111111";
				when "0101111001100111" => data <= "111111";
				when "0101111001101000" => data <= "111111";
				when "0101111001101111" => data <= "111111";
				when "0101111001110000" => data <= "111111";
				when "0101111001110100" => data <= "111111";
				when "0101111001110101" => data <= "111111";
				when "0101111001111010" => data <= "111111";
				when "0101111001111011" => data <= "111111";
				when "0101111010000001" => data <= "111111";
				when "0101111010000010" => data <= "111111";
				when "0101111100011110" => data <= "111111";
				when "0101111100011111" => data <= "111111";
				when "0101111100100111" => data <= "111111";
				when "0101111100101000" => data <= "111111";
				when "0101111100101101" => data <= "111111";
				when "0101111100101110" => data <= "111111";
				when "0101111100110001" => data <= "111111";
				when "0101111100110010" => data <= "111111";
				when "0101111101000000" => data <= "111111";
				when "0101111101000001" => data <= "111111";
				when "0101111101001011" => data <= "111111";
				when "0101111101001100" => data <= "111111";
				when "0101111101011100" => data <= "111111";
				when "0101111101011101" => data <= "111111";
				when "0101111101100010" => data <= "111111";
				when "0101111101100011" => data <= "111111";
				when "0101111101100111" => data <= "111111";
				when "0101111101101000" => data <= "111111";
				when "0101111101101111" => data <= "111111";
				when "0101111101110000" => data <= "111111";
				when "0101111101110100" => data <= "111111";
				when "0101111101110101" => data <= "111111";
				when "0101111101111010" => data <= "111111";
				when "0101111101111011" => data <= "111111";
				when "0101111110000001" => data <= "111111";
				when "0101111110000010" => data <= "111111";
				when "0110000000011110" => data <= "111111";
				when "0110000000011111" => data <= "111111";
				when "0110000000100111" => data <= "111111";
				when "0110000000101000" => data <= "111111";
				when "0110000000101101" => data <= "111111";
				when "0110000000101110" => data <= "111111";
				when "0110000000110001" => data <= "111111";
				when "0110000000110010" => data <= "111111";
				when "0110000000110011" => data <= "111111";
				when "0110000000110100" => data <= "111111";
				when "0110000000110101" => data <= "111111";
				when "0110000000110110" => data <= "111111";
				when "0110000000110111" => data <= "111111";
				when "0110000000111010" => data <= "111111";
				when "0110000000111011" => data <= "111111";
				when "0110000000111100" => data <= "111111";
				when "0110000000111101" => data <= "111111";
				when "0110000000111110" => data <= "111111";
				when "0110000000111111" => data <= "111111";
				when "0110000001000000" => data <= "111111";
				when "0110000001000001" => data <= "111111";
				when "0110000001000100" => data <= "111111";
				when "0110000001000101" => data <= "111111";
				when "0110000001000110" => data <= "111111";
				when "0110000001000111" => data <= "111111";
				when "0110000001001000" => data <= "111111";
				when "0110000001001001" => data <= "111111";
				when "0110000001001010" => data <= "111111";
				when "0110000001001011" => data <= "111111";
				when "0110000001001100" => data <= "111111";
				when "0110000001010101" => data <= "111111";
				when "0110000001010110" => data <= "111111";
				when "0110000001010111" => data <= "111111";
				when "0110000001011000" => data <= "111111";
				when "0110000001011001" => data <= "111111";
				when "0110000001011010" => data <= "111111";
				when "0110000001011011" => data <= "111111";
				when "0110000001011100" => data <= "111111";
				when "0110000001011101" => data <= "111111";
				when "0110000001100010" => data <= "111111";
				when "0110000001100011" => data <= "111111";
				when "0110000001100111" => data <= "111111";
				when "0110000001101000" => data <= "111111";
				when "0110000001101111" => data <= "111111";
				when "0110000001110000" => data <= "111111";
				when "0110000001110100" => data <= "111111";
				when "0110000001110101" => data <= "111111";
				when "0110000001111010" => data <= "111111";
				when "0110000001111011" => data <= "111111";
				when "0110000010000001" => data <= "111111";
				when "0110000010000010" => data <= "111111";
				when "0110000100011110" => data <= "111111";
				when "0110000100011111" => data <= "111111";
				when "0110000100100111" => data <= "111111";
				when "0110000100101000" => data <= "111111";
				when "0110000100101101" => data <= "111111";
				when "0110000100101110" => data <= "111111";
				when "0110000100110001" => data <= "111111";
				when "0110000100110010" => data <= "111111";
				when "0110000100110011" => data <= "111111";
				when "0110000100110100" => data <= "111111";
				when "0110000100110101" => data <= "111111";
				when "0110000100110110" => data <= "111111";
				when "0110000100110111" => data <= "111111";
				when "0110000100111010" => data <= "111111";
				when "0110000100111011" => data <= "111111";
				when "0110000100111100" => data <= "111111";
				when "0110000100111101" => data <= "111111";
				when "0110000100111110" => data <= "111111";
				when "0110000100111111" => data <= "111111";
				when "0110000101000100" => data <= "111111";
				when "0110000101000101" => data <= "111111";
				when "0110000101000110" => data <= "111111";
				when "0110000101000111" => data <= "111111";
				when "0110000101001000" => data <= "111111";
				when "0110000101001001" => data <= "111111";
				when "0110000101001010" => data <= "111111";
				when "0110000101010101" => data <= "111111";
				when "0110000101010110" => data <= "111111";
				when "0110000101010111" => data <= "111111";
				when "0110000101011000" => data <= "111111";
				when "0110000101011001" => data <= "111111";
				when "0110000101011010" => data <= "111111";
				when "0110000101011011" => data <= "111111";
				when "0110000101100010" => data <= "111111";
				when "0110000101100011" => data <= "111111";
				when "0110000101100111" => data <= "111111";
				when "0110000101101000" => data <= "111111";
				when "0110000101101111" => data <= "111111";
				when "0110000101110000" => data <= "111111";
				when "0110000101110100" => data <= "111111";
				when "0110000101110101" => data <= "111111";
				when "0110000101111010" => data <= "111111";
				when "0110000101111011" => data <= "111111";
				when "0110000110000001" => data <= "111111";
				when "0110000110000010" => data <= "111111";
				when others => data <= "000000";
			end case;
              		end if; 
              	end process; 
              end;
