library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity music is
	port(
		clk_in : in std_logic;
		sound : out std_logic;
		start : in std_logic;
		endsong : out std_logic
	);
end music;

architecture synth of music is 
	component clk_divider is
			port(
				clk_in : in std_logic;
				div_num : in integer;
				reset : in std_logic;
				clk_out : out std_logic
			);
	end component;
	
	component music_decoder is
		port(
			note_code : in std_logic_vector(3 downto 0);
			note_out : out integer
			);
	end component;
			

signal div : std_logic_vector(3 downto 0);
signal clk_sec : std_logic;
signal count : integer := 0;
signal reset_div : std_logic := '0';
signal temp : std_logic;
signal div_decoded : integer;

constant F4 : std_logic_vector(3 downto 0) := "0001";
constant G4 : std_logic_vector(3 downto 0) := "0010";
constant A4 : std_logic_vector(3 downto 0) := "0011";
constant C5 : std_logic_vector(3 downto 0) := "0100";
constant D5 : std_logic_vector(3 downto 0) := "0101";
constant E5 : std_logic_vector(3 downto 0) := "0110";
constant F5 : std_logic_vector(3 downto 0) := "0111";
constant G5 : std_logic_vector(3 downto 0) := "1000";
constant A5 : std_logic_vector(3 downto 0) := "1001";
constant C4 : std_logic_vector(3 downto 0) := "1010";
constant D4 : std_logic_vector(3 downto 0) := "1011";
constant B4f : std_logic_vector(3 downto 0) := "1100";
constant E4 : std_logic_vector(3 downto 0) := "1101";
	
begin

	sec_div : clk_divider
	port map(
		clk_in => clk_in,
		div_num => 131615,
		reset => '0',
		clk_out => clk_sec
	);
	
	music_div : clk_divider
	port map(
		clk_in => clk_in,
		div_num => div_decoded,
		reset => reset_div,
		clk_out => sound
	);
	
	decoder : music_decoder
	port map(
		note_code => div,
		note_out => div_decoded
	);
	
	process (clk_sec) is 
	begin 
		
		if rising_edge(clk_sec)then
			if (start = '0') then
				count <= 0;
				reset_div <= '1';
			else
			--endsong <= '0';
			if (count > -1 and count < 24) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 25) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 49) then
				reset_div <= '1';
			elsif (count = 50) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 74) then
				reset_div <= '1';
			elsif (count = 75) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 99) then
				reset_div <= '1';
			elsif (count = 100) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 124) then
				reset_div <= '1';
			elsif (count = 125) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 149) then
				reset_div <= '1';
			elsif (count = 150) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 174) then
				reset_div <= '1';
			elsif (count = 175) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 271) then
				reset_div <= '1';
			elsif (count = 272) then
				reset_div <= '1';
			elsif (count = 416) then
				reset_div <= '1';
			elsif (count = 417) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 441) then
				reset_div <= '1';
			elsif (count = 442) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 466) then
				reset_div <= '1';
			elsif (count = 467) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 491) then
				reset_div <= '1';
			elsif (count = 492) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 528) then
				reset_div <= '1';
			elsif (count = 529) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 565) then
				reset_div <= '1';
			elsif (count = 566) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 602) then
				reset_div <= '1';
			elsif (count = 603) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 615) then
				reset_div <= '1';
			elsif (count = 616) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 634) then
				reset_div <= '1';
			elsif (count = 635) then
				reset_div <= '1';
			elsif (count = 731) then
				reset_div <= '1';
			elsif (count = 732) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 756) then
				reset_div <= '1';
			elsif (count = 757) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 781) then
				reset_div <= '1';
			elsif (count = 782) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 806) then
				reset_div <= '1';
			elsif (count = 807) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 831) then
				reset_div <= '1';
			elsif (count = 832) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 856) then
				reset_div <= '1';
			elsif (count = 857) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 881) then
				reset_div <= '1';
			elsif (count = 882) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 906) then
				reset_div <= '1';
			elsif (count = 907) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 955) then
				reset_div <= '1';
			elsif (count = 956) then
				reset_div <= '1';
			elsif (count = 1124) then
				reset_div <= '1';
			elsif (count = 1125) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1149) then
				reset_div <= '1';
			elsif (count = 1150) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1174) then
				reset_div <= '1';
			elsif (count = 1175) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1199) then
				reset_div <= '1';
			elsif (count = 1200) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1224) then
				reset_div <= '1';
			elsif (count = 1225) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1249) then
				reset_div <= '1';
			elsif (count = 1250) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 1286) then
				reset_div <= '1';
			elsif (count = 1287) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1323) then
				reset_div <= '1';
			elsif (count = 1324) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1360) then
				reset_div <= '1';
			elsif (count = 1361) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 1373) then
				reset_div <= '1';
			elsif (count = 1374) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 1392) then
				reset_div <= '1';
			elsif (count = 1393) then
				reset_div <= '1';
			elsif (count = 1513) then
				reset_div <= '1';
			elsif (count = 1514) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 1538) then
				reset_div <= '1';
			elsif (count = 1539) then
				reset_div <= '0';
				div <= B4f;
			elsif (count = 1563) then
				reset_div <= '1';
			elsif (count = 1564) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 1588) then
				reset_div <= '1';
			elsif (count = 1589) then
				reset_div <= '0';
				div <= B4f;
			elsif (count = 1613) then
				reset_div <= '1';
			elsif (count = 1614) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 1638) then
				reset_div <= '1';
			elsif (count = 1639) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1663) then
				reset_div <= '1';
			elsif (count = 1664) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1688) then
				reset_div <= '1';
			elsif (count = 1689) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1701) then
				reset_div <= '1';
			elsif (count = 1702) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 1714) then
				reset_div <= '1';
			elsif (count = 1715) then
				reset_div <= '1';
			elsif (count = 1859) then
				reset_div <= '1';
			elsif (count = 1860) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1884) then
				reset_div <= '1';
			elsif (count = 1885) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1909) then
				reset_div <= '1';
			elsif (count = 1910) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 1934) then
				reset_div <= '1';
			elsif (count = 1935) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 1959) then
				reset_div <= '1';
			elsif (count = 1960) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 1996) then
				reset_div <= '1';
			elsif (count = 1997) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 2033) then
				reset_div <= '1';
			elsif (count = 2034) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2070) then
				reset_div <= '1';
			elsif (count = 2071) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 2083) then
				reset_div <= '1';
			elsif (count = 2084) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 2102) then
				reset_div <= '1';
			elsif (count = 2103) then
				reset_div <= '1';
			elsif (count = 2199) then
				reset_div <= '1';
			elsif (count = 2200) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 2224) then
				reset_div <= '1';
			elsif (count = 2225) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 2249) then
				reset_div <= '1';
			elsif (count = 2250) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 2274) then
				reset_div <= '1';
			elsif (count = 2275) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 2299) then
				reset_div <= '1';
			elsif (count = 2300) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 2324) then
				reset_div <= '1';
			elsif (count = 2325) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 2349) then
				reset_div <= '1';
			elsif (count = 2350) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2374) then
				reset_div <= '1';
			elsif (count = 2375) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2447) then
				reset_div <= '1';
			elsif (count = 2448) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 2460) then
				reset_div <= '1';
			elsif (count = 2461) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 2479) then
				reset_div <= '1';
			elsif (count = 2480) then
				reset_div <= '1';
			elsif (count = 2576) then
				reset_div <= '1';
			elsif (count = 2577) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2601) then
				reset_div <= '1';
			elsif (count = 2602) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 2626) then
				reset_div <= '1';
			elsif (count = 2627) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 2651) then
				reset_div <= '1';
			elsif (count = 2652) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 2676) then
				reset_div <= '1';
			elsif (count = 2677) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2701) then
				reset_div <= '1';
			elsif (count = 2702) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 2738) then
				reset_div <= '1';
			elsif (count = 2739) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 2775) then
				reset_div <= '1';
			elsif (count = 2776) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2812) then
				reset_div <= '1';
			elsif (count = 2813) then
				reset_div <= '0';
				div <= C4;
			elsif (count = 2825) then
				reset_div <= '1';
			elsif (count = 2826) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 2844) then
				reset_div <= '1';
			elsif (count = 2845) then
				reset_div <= '1';
			elsif (count = 2869) then
				reset_div <= '1';
			elsif (count = 2870) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2894) then
				reset_div <= '1';
			elsif (count = 2895) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 2931) then
				reset_div <= '1';
			elsif (count = 2932) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 2968) then
				reset_div <= '1';
			elsif (count = 2969) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 2993) then
				reset_div <= '1';
			elsif (count = 2994) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 3066) then
				reset_div <= '1';
			elsif (count = 3067) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3091) then
				reset_div <= '1';
			elsif (count = 3092) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 3128) then
				reset_div <= '1';
			elsif (count = 3129) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3165) then
				reset_div <= '1';
			elsif (count = 3166) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 3238) then
				reset_div <= '1';
			elsif (count = 3239) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 3263) then
				reset_div <= '1';
			elsif (count = 3264) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 3288) then
				reset_div <= '1';
			elsif (count = 3289) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 3325) then
				reset_div <= '1';
			elsif (count = 3326) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3362) then
				reset_div <= '1';
			elsif (count = 3363) then
				reset_div <= '0';
				div <= E4;
			elsif (count = 3435) then
				reset_div <= '1';
			elsif (count = 3436) then
				reset_div <= '1';
			elsif (count = 3460) then
				reset_div <= '1';
			elsif (count = 3461) then
				reset_div <= '0';
				div <= E4;
			elsif (count = 3485) then
				reset_div <= '1';
			elsif (count = 3486) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 3522) then
				reset_div <= '1';
			elsif (count = 3523) then
				reset_div <= '0';
				div <= E4;
			elsif (count = 3559) then
				reset_div <= '1';
			elsif (count = 3560) then
				reset_div <= '0';
				div <= D4;
			elsif (count = 3632) then
				reset_div <= '1';
			elsif (count = 3633) then
				reset_div <= '1';
			elsif (count = 3657) then
				reset_div <= '1';
			elsif (count = 3658) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 3682) then
				reset_div <= '1';
			elsif (count = 3683) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 3719) then
				reset_div <= '1';
			elsif (count = 3720) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 3756) then
				reset_div <= '1';
			elsif (count = 3757) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3781) then
				reset_div <= '1';
			elsif (count = 3782) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 3830) then
				reset_div <= '1';
			elsif (count = 3831) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 3855) then
				reset_div <= '1';
			elsif (count = 3856) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3880) then
				reset_div <= '1';
			elsif (count = 3881) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 3917) then
				reset_div <= '1';
			elsif (count = 3918) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 3954) then
				reset_div <= '1';
			elsif (count = 3955) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 4027) then
				reset_div <= '1';
			elsif (count = 4028) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 4052) then
				reset_div <= '1';
			elsif (count = 4053) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 4077) then
				reset_div <= '1';
			elsif (count = 4078) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 4102) then
				reset_div <= '1';
			elsif (count = 4103) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 4139) then
				reset_div <= '1';
			elsif (count = 4140) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 4176) then
				reset_div <= '1';
			elsif (count = 4177) then
				reset_div <= '0';
				div <= E4;
			elsif (count = 4249) then
				reset_div <= '1';
			elsif (count = 4250) then
				reset_div <= '1';
			elsif (count = 4394) then
				reset_div <= '1';
			elsif (count = 4395) then
				reset_div <= '0';
				div <= F4;
			elsif (count = 4419) then
				reset_div <= '1';
			elsif (count = 4420) then
				reset_div <= '0';
				div <= G4;
			elsif (count = 4444) then
				reset_div <= '1';
			elsif (count = 4445) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 4469) then
				reset_div <= '1';
			elsif (count = 4470) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 4494) then
				reset_div <= '1';
			elsif (count = 4495) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 4519) then
				reset_div <= '1';
			elsif (count = 4520) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 4544) then
				reset_div <= '1';
			elsif (count = 4545) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 4569) then
				reset_div <= '1';
			elsif (count = 4570) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 4594) then
				reset_div <= '1';
			elsif (count = 4595) then
				reset_div <= '0';
				div <= G5;
			elsif (count = 4631) then
				reset_div <= '1';
			elsif (count = 4632) then
				reset_div <= '0';
				div <= G5;
			elsif (count = 4668) then
				reset_div <= '1';
			elsif (count = 4669) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 4789) then
				reset_div <= '1';
			elsif (count = 4790) then
				reset_div <= '1';
			elsif (count = 4958) then
				reset_div <= '1';
			elsif (count = 4959) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 4971) then
				reset_div <= '1';
			elsif (count = 4972) then
				reset_div <= '0';
				div <= E5;
			elsif (count = 4984) then
				reset_div <= '1';
			elsif (count = 4985) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 5021) then
				reset_div <= '1';
			elsif (count = 5022) then
				reset_div <= '0';
				div <= A5;
			elsif (count = 5058) then
				reset_div <= '1';
			elsif (count = 5059) then
				reset_div <= '0';
				div <= E5;
			elsif (count = 5107) then
				reset_div <= '1';
			elsif (count = 5108) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 5132) then
				reset_div <= '1';
			elsif (count = 5133) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 5169) then
				reset_div <= '1';
			elsif (count = 5170) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 5194) then
				reset_div <= '1';
			elsif (count = 5195) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 5267) then
				reset_div <= '1';
			elsif (count = 5268) then
				reset_div <= '1';
			elsif (count = 5364) then
				reset_div <= '1';
			elsif (count = 5365) then
				reset_div <= '0';
				div <= G5;
			elsif (count = 5401) then
				reset_div <= '1';
			elsif (count = 5402) then
				reset_div <= '0';
				div <= G5;
			elsif (count = 5438) then
				reset_div <= '1';
			elsif (count = 5439) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 5559) then
				reset_div <= '1';
			elsif (count = 5560) then
				reset_div <= '1';
			elsif (count = 5728) then
				reset_div <= '1';
			elsif (count = 5729) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 5741) then
				reset_div <= '1';
			elsif (count = 5742) then
				reset_div <= '0';
				div <= E5;
			elsif (count = 5754) then
				reset_div <= '1';
			elsif (count = 5755) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 5791) then
				reset_div <= '1';
			elsif (count = 5792) then
				reset_div <= '0';
				div <= A5;
			elsif (count = 5828) then
				reset_div <= '1';
			elsif (count = 5829) then
				reset_div <= '0';
				div <= E5;
			elsif (count = 5877) then
				reset_div <= '1';
			elsif (count = 5878) then
				reset_div <= '0';
				div <= A4;
			elsif (count = 5902) then
				reset_div <= '1';
			elsif (count = 5903) then
				reset_div <= '0';
				div <= C5;
			elsif (count = 5939) then
				reset_div <= '1';
			elsif (count = 5940) then
				reset_div <= '0';
				div <= F5;
			elsif (count = 5976) then
				reset_div <= '1';
			elsif (count = 5977) then
				reset_div <= '0';
				div <= D5;
			elsif (count = 6049) then
				reset_div <= '1';
			elsif (count = 6050) then
				reset_div <= '1';
			--elsif (count = 6122) then
				--reset_div <= '1';
			--elsif (count = 6123) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 6135) then
				--reset_div <= '1';
			--elsif (count = 6136) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 6148) then
				--reset_div <= '1';
			--elsif (count = 6149) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 6185) then
				--reset_div <= '1';
			--elsif (count = 6186) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 6222) then
				--reset_div <= '1';
			--elsif (count = 6223) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 6271) then
				--reset_div <= '1';
			--elsif (count = 6272) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 6296) then
				--reset_div <= '1';
			--elsif (count = 6297) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 6333) then
				--reset_div <= '1';
			--elsif (count = 6334) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 6370) then
				--reset_div <= '1';
			--elsif (count = 6371) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 6443) then
				--reset_div <= '1';
			--elsif (count = 6444) then
				--reset_div <= '1';
			--elsif (count = 6516) then
				--reset_div <= '1';
			--elsif (count = 6517) then
				--reset_div <= '0';
				--div <= C4;
			--elsif (count = 6541) then
				--reset_div <= '1';
			--elsif (count = 6542) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 6566) then
				--reset_div <= '1';
			--elsif (count = 6567) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 6591) then
				--reset_div <= '1';
			--elsif (count = 6592) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 6616) then
				--reset_div <= '1';
			--elsif (count = 6617) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 6641) then
				--reset_div <= '1';
			--elsif (count = 6642) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 6666) then
				--reset_div <= '1';
			--elsif (count = 6667) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 6715) then
				--reset_div <= '1';
			--elsif (count = 6716) then
				--reset_div <= '1';
			--elsif (count = 6908) then
				--reset_div <= '1';
			--elsif (count = 6909) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 6933) then
				--reset_div <= '1';
			--elsif (count = 6934) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 6958) then
				--reset_div <= '1';
			--elsif (count = 6959) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 6983) then
				--reset_div <= '1';
			--elsif (count = 6984) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7008) then
				--reset_div <= '1';
			--elsif (count = 7009) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7045) then
				--reset_div <= '1';
			--elsif (count = 7046) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7082) then
				--reset_div <= '1';
			--elsif (count = 7083) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7119) then
				--reset_div <= '1';
			--elsif (count = 7120) then
				--reset_div <= '0';
				--div <= D4;
			--elsif (count = 7168) then
				--reset_div <= '1';
			--elsif (count = 7169) then
				--reset_div <= '1';
			--elsif (count = 7265) then
				--reset_div <= '1';
			--elsif (count = 7266) then
				--reset_div <= '0';
				--div <= C4;
			--elsif (count = 7290) then
				--reset_div <= '1';
			--elsif (count = 7291) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7315) then
				--reset_div <= '1';
			--elsif (count = 7316) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7340) then
				--reset_div <= '1';
			--elsif (count = 7341) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7365) then
				--reset_div <= '1';
			--elsif (count = 7366) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7390) then
				--reset_div <= '1';
			--elsif (count = 7391) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7415) then
				--reset_div <= '1';
			--elsif (count = 7416) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7440) then
				--reset_div <= '1';
			--elsif (count = 7441) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7489) then
				--reset_div <= '1';
			--elsif (count = 7490) then
				--reset_div <= '1';
			--elsif (count = 7658) then
				--reset_div <= '1';
			--elsif (count = 7659) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7683) then
				--reset_div <= '1';
			--elsif (count = 7684) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7708) then
				--reset_div <= '1';
			--elsif (count = 7709) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7733) then
				--reset_div <= '1';
			--elsif (count = 7734) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7758) then
				--reset_div <= '1';
			--elsif (count = 7759) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7783) then
				--reset_div <= '1';
			--elsif (count = 7784) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 7820) then
				--reset_div <= '1';
			--elsif (count = 7821) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 7857) then
				--reset_div <= '1';
			--elsif (count = 7858) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 7894) then
				--reset_div <= '1';
			--elsif (count = 7895) then
				--reset_div <= '0';
				--div <= D4;
			--elsif (count = 7943) then
				--reset_div <= '1';
			--elsif (count = 7944) then
				--reset_div <= '1';
			--elsif (count = 8040) then
				--reset_div <= '1';
			--elsif (count = 8041) then
				--reset_div <= '0';
				--div <= C4;
			--elsif (count = 8065) then
				--reset_div <= '1';
			--elsif (count = 8066) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 8090) then
				--reset_div <= '1';
			--elsif (count = 8091) then
				--reset_div <= '0';
				--div <= B4f;
			--elsif (count = 8115) then
				--reset_div <= '1';
			--elsif (count = 8116) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8140) then
				--reset_div <= '1';
			--elsif (count = 8141) then
				--reset_div <= '0';
				--div <= B4f;
			--elsif (count = 8165) then
				--reset_div <= '1';
			--elsif (count = 8166) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8190) then
				--reset_div <= '1';
			--elsif (count = 8191) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 8215) then
				--reset_div <= '1';
			--elsif (count = 8216) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 8312) then
				--reset_div <= '1';
			--elsif (count = 8313) then
				--reset_div <= '1';
			--elsif (count = 8457) then
				--reset_div <= '1';
			--elsif (count = 8458) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 8482) then
				--reset_div <= '1';
			--elsif (count = 8483) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 8507) then
				--reset_div <= '1';
			--elsif (count = 8508) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 8532) then
				--reset_div <= '1';
			--elsif (count = 8533) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 8557) then
				--reset_div <= '1';
			--elsif (count = 8558) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8594) then
				--reset_div <= '1';
			--elsif (count = 8595) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 8631) then
				--reset_div <= '1';
			--elsif (count = 8632) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 8668) then
				--reset_div <= '1';
			--elsif (count = 8669) then
				--reset_div <= '0';
				--div <= D4;
			--elsif (count = 8717) then
				--reset_div <= '1';
			--elsif (count = 8718) then
				--reset_div <= '1'; -- previous 3end 
			--elsif (count = 8814) then
				--reset_div <= '1';
			--elsif (count = 8815) then
				--reset_div <= '0';
				--div <= C4;
			--elsif (count = 8839) then
				--reset_div <= '1';
			--elsif (count = 8840) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8876) then
				--reset_div <= '1';
			--elsif (count = 8877) then
				--reset_div <= '0';
				--div <= B4f;
			--elsif (count = 8913) then
				--reset_div <= '1';
			--elsif (count = 8914) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8938) then
				--reset_div <= '1';
			--elsif (count = 8939) then
				--reset_div <= '0';
				--div <= B4f;
			--elsif (count = 8963) then
				--reset_div <= '1';
			--elsif (count = 8964) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 8988) then
				--reset_div <= '1';
			--elsif (count = 8989) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9013) then
				--reset_div <= '1';
			--elsif (count = 9014) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9110) then
				--reset_div <= '1';
			--elsif (count = 9111) then
				--reset_div <= '1';
			--elsif (count = 9231) then
				--reset_div <= '1';
			--elsif (count = 9232) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9256) then
				--reset_div <= '1';
			--elsif (count = 9257) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9281) then
				--reset_div <= '1';
			--elsif (count = 9282) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 9306) then
				--reset_div <= '1';
			--elsif (count = 9307) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 9331) then
				--reset_div <= '1';
			--elsif (count = 9332) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9356) then
				--reset_div <= '1';
			--elsif (count = 9357) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 9393) then
				--reset_div <= '1';
			--elsif (count = 9394) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 9430) then
				--reset_div <= '1';
			--elsif (count = 9431) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9467) then
				--reset_div <= '1';
			--elsif (count = 9468) then
				--reset_div <= '0';
				--div <= D4;
			--elsif (count = 9516) then
				--reset_div <= '1';
			--elsif (count = 9517) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9541) then
				--reset_div <= '1';
			--elsif (count = 9542) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 9578) then
				--reset_div <= '1';
			--elsif (count = 9579) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 9615) then
				--reset_div <= '1';
			--elsif (count = 9616) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 9640) then
				--reset_div <= '1';
			--elsif (count = 9641) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 9689) then
				--reset_div <= '1';
			--elsif (count = 9690) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 9714) then
				--reset_div <= '1';
			--elsif (count = 9715) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 9739) then
				--reset_div <= '1';
			--elsif (count = 9740) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 9776) then
				--reset_div <= '1';
			--elsif (count = 9777) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 9813) then
				--reset_div <= '1';
			--elsif (count = 9814) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 9886) then
				--reset_div <= '1';
			--elsif (count = 9887) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 9911) then
				--reset_div <= '1';
			--elsif (count = 9912) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 9936) then
				--reset_div <= '1';
			--elsif (count = 9937) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 9961) then
				--reset_div <= '1';
			--elsif (count = 9962) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 9998) then
				--reset_div <= '1';
			--elsif (count = 9999) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 10035) then
				--reset_div <= '1';
			--elsif (count = 10036) then
				--reset_div <= '0';
				--div <= E4;
			--elsif (count = 10108) then
				--reset_div <= '1';
			--elsif (count = 10109) then
				--reset_div <= '1';
			--elsif (count = 10253) then
				--reset_div <= '1';
			--elsif (count = 10254) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 10278) then
				--reset_div <= '1';
			--elsif (count = 10279) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 10303) then
				--reset_div <= '1';
			--elsif (count = 10304) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 10328) then
				--reset_div <= '1';
			--elsif (count = 10329) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 10353) then
				--reset_div <= '1';
			--elsif (count = 10354) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 10378) then
				--reset_div <= '1';
			--elsif (count = 10379) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 10403) then
				--reset_div <= '1';
			--elsif (count = 10404) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 10428) then
				--reset_div <= '1';
			--elsif (count = 10429) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 10453) then
				--reset_div <= '1';
			--elsif (count = 10454) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 10490) then
				--reset_div <= '1';
			--elsif (count = 10491) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 10527) then
				--reset_div <= '1';
			--elsif (count = 10528) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 10648) then
				--reset_div <= '1';
			--elsif (count = 10649) then
				--reset_div <= '1';
			--elsif (count = 10817) then
				--reset_div <= '1';
			--elsif (count = 10818) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 10830) then
				--reset_div <= '1';
			--elsif (count = 10831) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 10843) then
				--reset_div <= '1';
			--elsif (count = 10844) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 10880) then
				--reset_div <= '1';
			--elsif (count = 10881) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 10917) then
				--reset_div <= '1';
			--elsif (count = 10918) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 10966) then
				--reset_div <= '1';
			--elsif (count = 10967) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 10991) then
				--reset_div <= '1';
			--elsif (count = 10992) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 11028) then
				--reset_div <= '1';
			--elsif (count = 11029) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 11053) then
				--reset_div <= '1';
			--elsif (count = 11054) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 11126) then
				--reset_div <= '1';
			--elsif (count = 11127) then
				--reset_div <= '1';
			--elsif (count = 11223) then
				--reset_div <= '1';
			--elsif (count = 11224) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 11260) then
				--reset_div <= '1';
			--elsif (count = 11261) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 11297) then
				--reset_div <= '1';
			--elsif (count = 11298) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 11418) then
				--reset_div <= '1';
			--elsif (count = 11419) then
				--reset_div <= '1';
			--elsif (count = 11587) then
				--reset_div <= '1';
			--elsif (count = 11588) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 11600) then
				--reset_div <= '1';
			--elsif (count = 11601) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 11613) then
				--reset_div <= '1';
			--elsif (count = 11614) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 11650) then
				--reset_div <= '1';
			--elsif (count = 11651) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 11687) then
				--reset_div <= '1';
			--elsif (count = 11688) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 11736) then
				--reset_div <= '1';
			--elsif (count = 11737) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 11761) then
				--reset_div <= '1';
			--elsif (count = 11762) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 11798) then
				--reset_div <= '1';
			--elsif (count = 11799) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 11835) then
				--reset_div <= '1';
			--elsif (count = 11836) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 11908) then
				--reset_div <= '1';
			--elsif (count = 11909) then
				--reset_div <= '1';
			--elsif (count = 11981) then
				--reset_div <= '1';
			--elsif (count = 11982) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 11994) then
				--reset_div <= '1';
			--elsif (count = 11995) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 12007) then
				--reset_div <= '1';
			--elsif (count = 12008) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 12044) then
				--reset_div <= '1';
			--elsif (count = 12045) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 12081) then
				--reset_div <= '1';
			--elsif (count = 12082) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 12130) then
				--reset_div <= '1';
			--elsif (count = 12131) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 12155) then
				--reset_div <= '1';
			--elsif (count = 12156) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 12192) then
				--reset_div <= '1';
			--elsif (count = 12193) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 12229) then
				--reset_div <= '1';
			--elsif (count = 12230) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 12302) then
				--reset_div <= '1';
			--elsif (count = 12303) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12339) then
				--reset_div <= '1';
			--elsif (count = 12340) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12376) then
				--reset_div <= '1';
			--elsif (count = 12377) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12401) then
				--reset_div <= '1';
			--elsif (count = 12402) then
				--reset_div <= '1';
			--elsif (count = 12426) then
				--reset_div <= '1';
			--elsif (count = 12427) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 12451) then
				--reset_div <= '1';
			--elsif (count = 12452) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 12476) then
				--reset_div <= '1';
			--elsif (count = 12477) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 12501) then
				--reset_div <= '1';
			--elsif (count = 12502) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12538) then
				--reset_div <= '1';
			--elsif (count = 12539) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12575) then
				--reset_div <= '1';
			--elsif (count = 12576) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 12600) then
				--reset_div <= '1';
			--elsif (count = 12601) then
				--reset_div <= '1';
			--elsif (count = 13081) then
				--reset_div <= '1';
			--elsif (count = 13082) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13118) then
				--reset_div <= '1';
			--elsif (count = 13119) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13155) then
				--reset_div <= '1';
			--elsif (count = 13156) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13180) then
				--reset_div <= '1';
			--elsif (count = 13181) then
				--reset_div <= '1';
			--elsif (count = 13205) then
				--reset_div <= '1';
			--elsif (count = 13206) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 13230) then
				--reset_div <= '1';
			--elsif (count = 13231) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 13255) then
				--reset_div <= '1';
			--elsif (count = 13256) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 13280) then
				--reset_div <= '1';
			--elsif (count = 13281) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13317) then
				--reset_div <= '1';
			--elsif (count = 13318) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13354) then
				--reset_div <= '1';
			--elsif (count = 13355) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13379) then
				--reset_div <= '1';
			--elsif (count = 13380) then
				--reset_div <= '1';
			--elsif (count = 13740) then
				--reset_div <= '1';
			--elsif (count = 13741) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13765) then
				--reset_div <= '1';
			--elsif (count = 13766) then
				--reset_div <= '0';
				--div <= F4;
			--elsif (count = 13802) then
				--reset_div <= '1';
			--elsif (count = 13803) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 13839) then
				--reset_div <= '1';
			--elsif (count = 13840) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 13864) then
				--reset_div <= '1';
			--elsif (count = 13865) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 13913) then
				--reset_div <= '1';
			--elsif (count = 13914) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 13938) then
				--reset_div <= '1';
			--elsif (count = 13939) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 13963) then
				--reset_div <= '1';
			--elsif (count = 13964) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 14000) then
				--reset_div <= '1';
			--elsif (count = 14001) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 14037) then
				--reset_div <= '1';
			--elsif (count = 14038) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 14110) then
				--reset_div <= '1';
			--elsif (count = 14111) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 14135) then
				--reset_div <= '1';
			--elsif (count = 14136) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 14160) then
				--reset_div <= '1';
			--elsif (count = 14161) then
				--reset_div <= '0';
				--div <= G4;
			--elsif (count = 14185) then
				--reset_div <= '1';
			--elsif (count = 14186) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 14222) then
				--reset_div <= '1';
			--elsif (count = 14223) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 14259) then
				--reset_div <= '1';
			--elsif (count = 14260) then
				--reset_div <= '0';
				--div <= E4;
			--elsif (count = 14332) then
				--reset_div <= '1';
			--elsif (count = 14333) then
				--reset_div <= '1';
			--elsif (count = 14477) then
				--reset_div <= '1';
			--elsif (count = 14478) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 14514) then
				--reset_div <= '1';
			--elsif (count = 14515) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 14551) then
				--reset_div <= '1';
			--elsif (count = 14552) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 14672) then
				--reset_div <= '1';
			--elsif (count = 14673) then
				--reset_div <= '1';
			--elsif (count = 14841) then
				--reset_div <= '1';
			--elsif (count = 14842) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 14854) then
				--reset_div <= '1';
			--elsif (count = 14855) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 14867) then
				--reset_div <= '1';
			--elsif (count = 14868) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 14904) then
				--reset_div <= '1';
			--elsif (count = 14905) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 14941) then
				--reset_div <= '1';
			--elsif (count = 14942) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 14990) then
				--reset_div <= '1';
			--elsif (count = 14991) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 15015) then
				--reset_div <= '1';
			--elsif (count = 15016) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 15052) then
				--reset_div <= '1';
			--elsif (count = 15053) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 15077) then
				--reset_div <= '1';
			--elsif (count = 15078) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 15150) then
				--reset_div <= '1';
			--elsif (count = 15151) then
				--reset_div <= '1';
			--elsif (count = 15247) then
				--reset_div <= '1';
			--elsif (count = 15248) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 15284) then
				--reset_div <= '1';
			--elsif (count = 15285) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 15321) then
				--reset_div <= '1';
			--elsif (count = 15322) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 15442) then
				--reset_div <= '1';
			--elsif (count = 15443) then
				--reset_div <= '1';
			--elsif (count = 15611) then
				--reset_div <= '1';
			--elsif (count = 15612) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 15624) then
				--reset_div <= '1';
			--elsif (count = 15625) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 15637) then
				--reset_div <= '1';
			--elsif (count = 15638) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 15674) then
				--reset_div <= '1';
			--elsif (count = 15675) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 15711) then
				--reset_div <= '1';
			--elsif (count = 15712) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 15760) then
				--reset_div <= '1';
			--elsif (count = 15761) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 15785) then
				--reset_div <= '1';
			--elsif (count = 15786) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 15822) then
				--reset_div <= '1';
			--elsif (count = 15823) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 15847) then
				--reset_div <= '1';
			--elsif (count = 15848) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 15920) then
				--reset_div <= '1';
			--elsif (count = 15921) then
				--reset_div <= '1';
			--elsif (count = 16017) then
				--reset_div <= '1';
			--elsif (count = 16018) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 16054) then
				--reset_div <= '1';
			--elsif (count = 16055) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 16091) then
				--reset_div <= '1';
			--elsif (count = 16092) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 16212) then
				--reset_div <= '1';
			--elsif (count = 16213) then
				--reset_div <= '1';
			--elsif (count = 16381) then
				--reset_div <= '1';
			--elsif (count = 16382) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 16394) then
				--reset_div <= '1';
			--elsif (count = 16395) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 16407) then
				--reset_div <= '1';
			--elsif (count = 16408) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 16444) then
				--reset_div <= '1';
			--elsif (count = 16445) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 16481) then
				--reset_div <= '1';
			--elsif (count = 16482) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 16530) then
				--reset_div <= '1';
			--elsif (count = 16531) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 16555) then
				--reset_div <= '1';
			--elsif (count = 16556) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 16592) then
				--reset_div <= '1';
			--elsif (count = 16593) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 16617) then
				--reset_div <= '1';
			--elsif (count = 16618) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 16690) then
				--reset_div <= '1';
			--elsif (count = 16691) then
				--reset_div <= '1';
			--elsif (count = 16787) then
				--reset_div <= '1';
			--elsif (count = 16788) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 16824) then
				--reset_div <= '1';
			--elsif (count = 16825) then
				--reset_div <= '0';
				--div <= G5;
			--elsif (count = 16861) then
				--reset_div <= '1';
			--elsif (count = 16862) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 16982) then
				--reset_div <= '1';
			--elsif (count = 16983) then
				--reset_div <= '1';
			--elsif (count = 17151) then
				--reset_div <= '1';
			--elsif (count = 17152) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 17164) then
				--reset_div <= '1';
			--elsif (count = 17165) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 17177) then
				--reset_div <= '1';
			--elsif (count = 17178) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 17214) then
				--reset_div <= '1';
			--elsif (count = 17215) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 17251) then
				--reset_div <= '1';
			--elsif (count = 17252) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 17300) then
				--reset_div <= '1';
			--elsif (count = 17301) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 17325) then
				--reset_div <= '1';
			--elsif (count = 17326) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 17362) then
				--reset_div <= '1';
			--elsif (count = 17363) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 17399) then
				--reset_div <= '1';
			--elsif (count = 17400) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 17472) then
				--reset_div <= '1';
			--elsif (count = 17473) then
				--reset_div <= '1';
			--elsif (count = 17545) then
				--reset_div <= '1';
			--elsif (count = 17546) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 17558) then
				--reset_div <= '1';
			--elsif (count = 17559) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 17571) then
				--reset_div <= '1';
			--elsif (count = 17572) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 17608) then
				--reset_div <= '1';
			--elsif (count = 17609) then
				--reset_div <= '0';
				--div <= A5;
			--elsif (count = 17645) then
				--reset_div <= '1';
			--elsif (count = 17646) then
				--reset_div <= '0';
				--div <= E5;
			--elsif (count = 17694) then
				--reset_div <= '1';
			--elsif (count = 17695) then
				--reset_div <= '0';
				--div <= A4;
			--elsif (count = 17719) then
				--reset_div <= '1';
			--elsif (count = 17720) then
				--reset_div <= '0';
				--div <= C5;
			--elsif (count = 17756) then
				--reset_div <= '1';
			--elsif (count = 17757) then
				--reset_div <= '0';
				--div <= F5;
			--elsif (count = 17793) then
				--reset_div <= '1';
			--elsif (count = 17794) then
				--reset_div <= '0';
				--div <= D5;
			--elsif (count = 17866) then
				--reset_div <= '1';
			end if;
			count <= count + 1;
			end if;
		end if;
	end process;
	endsong <= '1' when count = 6050 else '0';
end;
	
		
	
	
	
	