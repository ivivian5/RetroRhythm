library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity rom is 
 	port(
		outglobal_o : in std_logic;
		addr_x : in std_logic_vector(6 downto 0);
		addr_y : in std_logic_vector(6 downto 0);
		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
	);
end;

architecture sim of rom is
signal addr : std_logic_vector(13 downto 0);

begin
	addr (13 downto 7) <= addr_y;
	addr (6 downto 0) <= addr_x;
	process(outglobal_o) begin
		if rising_edge(outglobal_o) then
			case addr is
				when "00001010010101" => data <= "111111";
				when "00001010010110" => data <= "111111";
				when "00001010010111" => data <= "111111";
				when "00001010011000" => data <= "111111";
				when "00001010011110" => data <= "111111";
				when "00001010011111" => data <= "111111";
				when "00001010100000" => data <= "111111";
				when "00001010100001" => data <= "111111";
				when "00001010100010" => data <= "111111";
				when "00001010100111" => data <= "111111";
				when "00001010101000" => data <= "111111";
				when "00001010101001" => data <= "111111";
				when "00001010101010" => data <= "111111";
				when "00001010101011" => data <= "111111";
				when "00001010110000" => data <= "111111";
				when "00001010110001" => data <= "111111";
				when "00001010110010" => data <= "111111";
				when "00001010110011" => data <= "111111";
				when "00001010111010" => data <= "111111";
				when "00001010111011" => data <= "111111";
				when "00001010111100" => data <= "111111";
				when "00001010111101" => data <= "111111";
				when "00001100010100" => data <= "111111";
				when "00001100010101" => data <= "010011";
				when "00001100010110" => data <= "010011";
				when "00001100010111" => data <= "010011";
				when "00001100011000" => data <= "010011";
				when "00001100011001" => data <= "111111";
				when "00001100011101" => data <= "111111";
				when "00001100011110" => data <= "010011";
				when "00001100011111" => data <= "010011";
				when "00001100100000" => data <= "010011";
				when "00001100100001" => data <= "010011";
				when "00001100100010" => data <= "010011";
				when "00001100100011" => data <= "111111";
				when "00001100100110" => data <= "111111";
				when "00001100100111" => data <= "010011";
				when "00001100101000" => data <= "010011";
				when "00001100101001" => data <= "010011";
				when "00001100101010" => data <= "010011";
				when "00001100101011" => data <= "010011";
				when "00001100101100" => data <= "111111";
				when "00001100101111" => data <= "111111";
				when "00001100110000" => data <= "010011";
				when "00001100110001" => data <= "010011";
				when "00001100110010" => data <= "010011";
				when "00001100110011" => data <= "010011";
				when "00001100110100" => data <= "111111";
				when "00001100111001" => data <= "111111";
				when "00001100111010" => data <= "010011";
				when "00001100111011" => data <= "010011";
				when "00001100111100" => data <= "010011";
				when "00001100111101" => data <= "010011";
				when "00001100111110" => data <= "111111";
				when "00001110010100" => data <= "111111";
				when "00001110010101" => data <= "010011";
				when "00001110010110" => data <= "111111";
				when "00001110010111" => data <= "111111";
				when "00001110011000" => data <= "111111";
				when "00001110011001" => data <= "010011";
				when "00001110011010" => data <= "111111";
				when "00001110011101" => data <= "111111";
				when "00001110011110" => data <= "010011";
				when "00001110011111" => data <= "111111";
				when "00001110100000" => data <= "111111";
				when "00001110100001" => data <= "111111";
				when "00001110100010" => data <= "111111";
				when "00001110100111" => data <= "111111";
				when "00001110101000" => data <= "111111";
				when "00001110101001" => data <= "010011";
				when "00001110101010" => data <= "111111";
				when "00001110101011" => data <= "111111";
				when "00001110101111" => data <= "111111";
				when "00001110110000" => data <= "010011";
				when "00001110110001" => data <= "111111";
				when "00001110110010" => data <= "111111";
				when "00001110110011" => data <= "111111";
				when "00001110110100" => data <= "010011";
				when "00001110110101" => data <= "111111";
				when "00001110111000" => data <= "111111";
				when "00001110111001" => data <= "010011";
				when "00001110111010" => data <= "111111";
				when "00001110111011" => data <= "111111";
				when "00001110111100" => data <= "111111";
				when "00001110111101" => data <= "111111";
				when "00001110111110" => data <= "010011";
				when "00001110111111" => data <= "111111";
				when "00010000010100" => data <= "111111";
				when "00010000010101" => data <= "010010";
				when "00010000010110" => data <= "111111";
				when "00010000010111" => data <= "111111";
				when "00010000011000" => data <= "111111";
				when "00010000011001" => data <= "010010";
				when "00010000011010" => data <= "111111";
				when "00010000011101" => data <= "111111";
				when "00010000011110" => data <= "010010";
				when "00010000011111" => data <= "111111";
				when "00010000100000" => data <= "111111";
				when "00010000101000" => data <= "111111";
				when "00010000101001" => data <= "010010";
				when "00010000101010" => data <= "111111";
				when "00010000101111" => data <= "111111";
				when "00010000110000" => data <= "010010";
				when "00010000110001" => data <= "111111";
				when "00010000110011" => data <= "111111";
				when "00010000110100" => data <= "010010";
				when "00010000110101" => data <= "111111";
				when "00010000111000" => data <= "111111";
				when "00010000111001" => data <= "010010";
				when "00010000111010" => data <= "111111";
				when "00010000111101" => data <= "111111";
				when "00010000111110" => data <= "010010";
				when "00010000111111" => data <= "111111";
				when "00010010010100" => data <= "111111";
				when "00010010010101" => data <= "010010";
				when "00010010010110" => data <= "010010";
				when "00010010010111" => data <= "010010";
				when "00010010011000" => data <= "010010";
				when "00010010011001" => data <= "010010";
				when "00010010011010" => data <= "111111";
				when "00010010011101" => data <= "111111";
				when "00010010011110" => data <= "010010";
				when "00010010011111" => data <= "010010";
				when "00010010100000" => data <= "010010";
				when "00010010100001" => data <= "111111";
				when "00010010101000" => data <= "111111";
				when "00010010101001" => data <= "010010";
				when "00010010101010" => data <= "111111";
				when "00010010101111" => data <= "111111";
				when "00010010110000" => data <= "010010";
				when "00010010110001" => data <= "111111";
				when "00010010110010" => data <= "111111";
				when "00010010110011" => data <= "111111";
				when "00010010110100" => data <= "010010";
				when "00010010110101" => data <= "111111";
				when "00010010111000" => data <= "111111";
				when "00010010111001" => data <= "010010";
				when "00010010111010" => data <= "111111";
				when "00010010111101" => data <= "111111";
				when "00010010111110" => data <= "010010";
				when "00010010111111" => data <= "111111";
				when "00010100010100" => data <= "111111";
				when "00010100010101" => data <= "100010";
				when "00010100010110" => data <= "100010";
				when "00010100010111" => data <= "100010";
				when "00010100011000" => data <= "100010";
				when "00010100011001" => data <= "111111";
				when "00010100011101" => data <= "111111";
				when "00010100011110" => data <= "100010";
				when "00010100011111" => data <= "111111";
				when "00010100100000" => data <= "111111";
				when "00010100101000" => data <= "111111";
				when "00010100101001" => data <= "100010";
				when "00010100101010" => data <= "111111";
				when "00010100101111" => data <= "111111";
				when "00010100110000" => data <= "100010";
				when "00010100110001" => data <= "100010";
				when "00010100110010" => data <= "100010";
				when "00010100110011" => data <= "100010";
				when "00010100110100" => data <= "111111";
				when "00010100111000" => data <= "111111";
				when "00010100111001" => data <= "100010";
				when "00010100111010" => data <= "111111";
				when "00010100111101" => data <= "111111";
				when "00010100111110" => data <= "100010";
				when "00010100111111" => data <= "111111";
				when "00010110010100" => data <= "111111";
				when "00010110010101" => data <= "100010";
				when "00010110010110" => data <= "111111";
				when "00010110010111" => data <= "111111";
				when "00010110011000" => data <= "111111";
				when "00010110011001" => data <= "100010";
				when "00010110011010" => data <= "111111";
				when "00010110011101" => data <= "111111";
				when "00010110011110" => data <= "100010";
				when "00010110011111" => data <= "111111";
				when "00010110101000" => data <= "111111";
				when "00010110101001" => data <= "100010";
				when "00010110101010" => data <= "111111";
				when "00010110101111" => data <= "111111";
				when "00010110110000" => data <= "100010";
				when "00010110110001" => data <= "111111";
				when "00010110110010" => data <= "111111";
				when "00010110110011" => data <= "111111";
				when "00010110110100" => data <= "100010";
				when "00010110110101" => data <= "111111";
				when "00010110111000" => data <= "111111";
				when "00010110111001" => data <= "100010";
				when "00010110111010" => data <= "111111";
				when "00010110111101" => data <= "111111";
				when "00010110111110" => data <= "100010";
				when "00010110111111" => data <= "111111";
				when "00011000010100" => data <= "111111";
				when "00011000010101" => data <= "110010";
				when "00011000010110" => data <= "111111";
				when "00011000011000" => data <= "111111";
				when "00011000011001" => data <= "110010";
				when "00011000011010" => data <= "111111";
				when "00011000011101" => data <= "111111";
				when "00011000011110" => data <= "110010";
				when "00011000011111" => data <= "111111";
				when "00011000100000" => data <= "111111";
				when "00011000100001" => data <= "111111";
				when "00011000100010" => data <= "111111";
				when "00011000101000" => data <= "111111";
				when "00011000101001" => data <= "110010";
				when "00011000101010" => data <= "111111";
				when "00011000101111" => data <= "111111";
				when "00011000110000" => data <= "110010";
				when "00011000110001" => data <= "111111";
				when "00011000110011" => data <= "111111";
				when "00011000110100" => data <= "110010";
				when "00011000110101" => data <= "111111";
				when "00011000111000" => data <= "111111";
				when "00011000111001" => data <= "110010";
				when "00011000111010" => data <= "111111";
				when "00011000111011" => data <= "111111";
				when "00011000111100" => data <= "111111";
				when "00011000111101" => data <= "111111";
				when "00011000111110" => data <= "110010";
				when "00011000111111" => data <= "111111";
				when "00011010010100" => data <= "111111";
				when "00011010010101" => data <= "110010";
				when "00011010010110" => data <= "111111";
				when "00011010011000" => data <= "111111";
				when "00011010011001" => data <= "110010";
				when "00011010011010" => data <= "111111";
				when "00011010011101" => data <= "111111";
				when "00011010011110" => data <= "110010";
				when "00011010011111" => data <= "110010";
				when "00011010100000" => data <= "110010";
				when "00011010100001" => data <= "110010";
				when "00011010100010" => data <= "110010";
				when "00011010100011" => data <= "111111";
				when "00011010101000" => data <= "111111";
				when "00011010101001" => data <= "110010";
				when "00011010101010" => data <= "111111";
				when "00011010101111" => data <= "111111";
				when "00011010110000" => data <= "110010";
				when "00011010110001" => data <= "111111";
				when "00011010110011" => data <= "111111";
				when "00011010110100" => data <= "110010";
				when "00011010110101" => data <= "111111";
				when "00011010111001" => data <= "111111";
				when "00011010111010" => data <= "110010";
				when "00011010111011" => data <= "110010";
				when "00011010111100" => data <= "110010";
				when "00011010111101" => data <= "110010";
				when "00011010111110" => data <= "111111";
				when "00011100010101" => data <= "111111";
				when "00011100011001" => data <= "111111";
				when "00011100011110" => data <= "111111";
				when "00011100011111" => data <= "111111";
				when "00011100100000" => data <= "111111";
				when "00011100100001" => data <= "111111";
				when "00011100100010" => data <= "111111";
				when "00011100101001" => data <= "111111";
				when "00011100110000" => data <= "111111";
				when "00011100110100" => data <= "111111";
				when "00011100111010" => data <= "111111";
				when "00011100111011" => data <= "111111";
				when "00011100111100" => data <= "111111";
				when "00011100111101" => data <= "111111";
				when "00100010001110" => data <= "111111";
				when "00100010001111" => data <= "111111";
				when "00100010010000" => data <= "111111";
				when "00100010010001" => data <= "111111";
				when "00100010010110" => data <= "111111";
				when "00100010011010" => data <= "111111";
				when "00100010011110" => data <= "111111";
				when "00100010100010" => data <= "111111";
				when "00100010100110" => data <= "111111";
				when "00100010100111" => data <= "111111";
				when "00100010101000" => data <= "111111";
				when "00100010101001" => data <= "111111";
				when "00100010101010" => data <= "111111";
				when "00100010101110" => data <= "111111";
				when "00100010110010" => data <= "111111";
				when "00100010110110" => data <= "111111";
				when "00100010111010" => data <= "111111";
				when "00100010111110" => data <= "111111";
				when "00100011000010" => data <= "111111";
				when "00100100001101" => data <= "111111";
				when "00100100001110" => data <= "010011";
				when "00100100001111" => data <= "010011";
				when "00100100010000" => data <= "010011";
				when "00100100010001" => data <= "010011";
				when "00100100010010" => data <= "111111";
				when "00100100010101" => data <= "111111";
				when "00100100010110" => data <= "010011";
				when "00100100010111" => data <= "111111";
				when "00100100011001" => data <= "111111";
				when "00100100011010" => data <= "010011";
				when "00100100011011" => data <= "111111";
				when "00100100011101" => data <= "111111";
				when "00100100011110" => data <= "010011";
				when "00100100011111" => data <= "111111";
				when "00100100100001" => data <= "111111";
				when "00100100100010" => data <= "010011";
				when "00100100100011" => data <= "111111";
				when "00100100100101" => data <= "111111";
				when "00100100100110" => data <= "010011";
				when "00100100100111" => data <= "010011";
				when "00100100101000" => data <= "010011";
				when "00100100101001" => data <= "010011";
				when "00100100101010" => data <= "010011";
				when "00100100101011" => data <= "111111";
				when "00100100101101" => data <= "111111";
				when "00100100101110" => data <= "010011";
				when "00100100101111" => data <= "111111";
				when "00100100110001" => data <= "111111";
				when "00100100110010" => data <= "010011";
				when "00100100110011" => data <= "111111";
				when "00100100110101" => data <= "111111";
				when "00100100110110" => data <= "010011";
				when "00100100110111" => data <= "111111";
				when "00100100111001" => data <= "111111";
				when "00100100111010" => data <= "010011";
				when "00100100111011" => data <= "111111";
				when "00100100111101" => data <= "111111";
				when "00100100111110" => data <= "010011";
				when "00100100111111" => data <= "111111";
				when "00100101000001" => data <= "111111";
				when "00100101000010" => data <= "010011";
				when "00100101000011" => data <= "111111";
				when "00100110001101" => data <= "111111";
				when "00100110001110" => data <= "010011";
				when "00100110001111" => data <= "111111";
				when "00100110010000" => data <= "111111";
				when "00100110010001" => data <= "111111";
				when "00100110010010" => data <= "010011";
				when "00100110010011" => data <= "111111";
				when "00100110010101" => data <= "111111";
				when "00100110010110" => data <= "010011";
				when "00100110010111" => data <= "111111";
				when "00100110011001" => data <= "111111";
				when "00100110011010" => data <= "010011";
				when "00100110011011" => data <= "111111";
				when "00100110011101" => data <= "111111";
				when "00100110011110" => data <= "010011";
				when "00100110011111" => data <= "111111";
				when "00100110100001" => data <= "111111";
				when "00100110100010" => data <= "010011";
				when "00100110100011" => data <= "111111";
				when "00100110100110" => data <= "111111";
				when "00100110100111" => data <= "111111";
				when "00100110101000" => data <= "010011";
				when "00100110101001" => data <= "111111";
				when "00100110101010" => data <= "111111";
				when "00100110101101" => data <= "111111";
				when "00100110101110" => data <= "010011";
				when "00100110101111" => data <= "111111";
				when "00100110110001" => data <= "111111";
				when "00100110110010" => data <= "010011";
				when "00100110110011" => data <= "111111";
				when "00100110110101" => data <= "111111";
				when "00100110110110" => data <= "010011";
				when "00100110110111" => data <= "111111";
				when "00100110111001" => data <= "111111";
				when "00100110111010" => data <= "010011";
				when "00100110111011" => data <= "111111";
				when "00100110111101" => data <= "111111";
				when "00100110111110" => data <= "010011";
				when "00100110111111" => data <= "010011";
				when "00100111000000" => data <= "111111";
				when "00100111000001" => data <= "010011";
				when "00100111000010" => data <= "010011";
				when "00100111000011" => data <= "111111";
				when "00101000001101" => data <= "111111";
				when "00101000001110" => data <= "010010";
				when "00101000001111" => data <= "111111";
				when "00101000010000" => data <= "111111";
				when "00101000010001" => data <= "111111";
				when "00101000010010" => data <= "010010";
				when "00101000010011" => data <= "111111";
				when "00101000010101" => data <= "111111";
				when "00101000010110" => data <= "010010";
				when "00101000010111" => data <= "111111";
				when "00101000011000" => data <= "111111";
				when "00101000011001" => data <= "111111";
				when "00101000011010" => data <= "010010";
				when "00101000011011" => data <= "111111";
				when "00101000011101" => data <= "111111";
				when "00101000011110" => data <= "010010";
				when "00101000011111" => data <= "010010";
				when "00101000100000" => data <= "111111";
				when "00101000100001" => data <= "010010";
				when "00101000100010" => data <= "010010";
				when "00101000100011" => data <= "111111";
				when "00101000100111" => data <= "111111";
				when "00101000101000" => data <= "010010";
				when "00101000101001" => data <= "111111";
				when "00101000101101" => data <= "111111";
				when "00101000101110" => data <= "010010";
				when "00101000101111" => data <= "111111";
				when "00101000110000" => data <= "111111";
				when "00101000110001" => data <= "111111";
				when "00101000110010" => data <= "010010";
				when "00101000110011" => data <= "111111";
				when "00101000110101" => data <= "111111";
				when "00101000110110" => data <= "010010";
				when "00101000110111" => data <= "010010";
				when "00101000111000" => data <= "111111";
				when "00101000111001" => data <= "010010";
				when "00101000111010" => data <= "010010";
				when "00101000111011" => data <= "111111";
				when "00101000111101" => data <= "111111";
				when "00101000111110" => data <= "010010";
				when "00101000111111" => data <= "111111";
				when "00101001000000" => data <= "010010";
				when "00101001000001" => data <= "111111";
				when "00101001000010" => data <= "010010";
				when "00101001000011" => data <= "111111";
				when "00101010001101" => data <= "111111";
				when "00101010001110" => data <= "010010";
				when "00101010001111" => data <= "010010";
				when "00101010010000" => data <= "010010";
				when "00101010010001" => data <= "010010";
				when "00101010010010" => data <= "010010";
				when "00101010010011" => data <= "111111";
				when "00101010010101" => data <= "111111";
				when "00101010010110" => data <= "010010";
				when "00101010010111" => data <= "010010";
				when "00101010011000" => data <= "010010";
				when "00101010011001" => data <= "010010";
				when "00101010011010" => data <= "010010";
				when "00101010011011" => data <= "111111";
				when "00101010011110" => data <= "111111";
				when "00101010011111" => data <= "010010";
				when "00101010100000" => data <= "010010";
				when "00101010100001" => data <= "010010";
				when "00101010100010" => data <= "111111";
				when "00101010100111" => data <= "111111";
				when "00101010101000" => data <= "010010";
				when "00101010101001" => data <= "111111";
				when "00101010101101" => data <= "111111";
				when "00101010101110" => data <= "010010";
				when "00101010101111" => data <= "010010";
				when "00101010110000" => data <= "010010";
				when "00101010110001" => data <= "010010";
				when "00101010110010" => data <= "010010";
				when "00101010110011" => data <= "111111";
				when "00101010110110" => data <= "111111";
				when "00101010110111" => data <= "010010";
				when "00101010111000" => data <= "010010";
				when "00101010111001" => data <= "010010";
				when "00101010111010" => data <= "111111";
				when "00101010111101" => data <= "111111";
				when "00101010111110" => data <= "010010";
				when "00101010111111" => data <= "111111";
				when "00101011000000" => data <= "111111";
				when "00101011000001" => data <= "111111";
				when "00101011000010" => data <= "010010";
				when "00101011000011" => data <= "111111";
				when "00101100001101" => data <= "111111";
				when "00101100001110" => data <= "100010";
				when "00101100001111" => data <= "100010";
				when "00101100010000" => data <= "100010";
				when "00101100010001" => data <= "100010";
				when "00101100010010" => data <= "111111";
				when "00101100010101" => data <= "111111";
				when "00101100010110" => data <= "100010";
				when "00101100010111" => data <= "111111";
				when "00101100011000" => data <= "111111";
				when "00101100011001" => data <= "111111";
				when "00101100011010" => data <= "100010";
				when "00101100011011" => data <= "111111";
				when "00101100011111" => data <= "111111";
				when "00101100100000" => data <= "100010";
				when "00101100100001" => data <= "111111";
				when "00101100100111" => data <= "111111";
				when "00101100101000" => data <= "100010";
				when "00101100101001" => data <= "111111";
				when "00101100101101" => data <= "111111";
				when "00101100101110" => data <= "100010";
				when "00101100101111" => data <= "111111";
				when "00101100110000" => data <= "111111";
				when "00101100110001" => data <= "111111";
				when "00101100110010" => data <= "100010";
				when "00101100110011" => data <= "111111";
				when "00101100110111" => data <= "111111";
				when "00101100111000" => data <= "100010";
				when "00101100111001" => data <= "111111";
				when "00101100111101" => data <= "111111";
				when "00101100111110" => data <= "100010";
				when "00101100111111" => data <= "111111";
				when "00101101000001" => data <= "111111";
				when "00101101000010" => data <= "100010";
				when "00101101000011" => data <= "111111";
				when "00101110001101" => data <= "111111";
				when "00101110001110" => data <= "100010";
				when "00101110001111" => data <= "111111";
				when "00101110010000" => data <= "111111";
				when "00101110010001" => data <= "111111";
				when "00101110010010" => data <= "100010";
				when "00101110010011" => data <= "111111";
				when "00101110010101" => data <= "111111";
				when "00101110010110" => data <= "100010";
				when "00101110010111" => data <= "111111";
				when "00101110011001" => data <= "111111";
				when "00101110011010" => data <= "100010";
				when "00101110011011" => data <= "111111";
				when "00101110011111" => data <= "111111";
				when "00101110100000" => data <= "100010";
				when "00101110100001" => data <= "111111";
				when "00101110100111" => data <= "111111";
				when "00101110101000" => data <= "100010";
				when "00101110101001" => data <= "111111";
				when "00101110101101" => data <= "111111";
				when "00101110101110" => data <= "100010";
				when "00101110101111" => data <= "111111";
				when "00101110110001" => data <= "111111";
				when "00101110110010" => data <= "100010";
				when "00101110110011" => data <= "111111";
				when "00101110110111" => data <= "111111";
				when "00101110111000" => data <= "100010";
				when "00101110111001" => data <= "111111";
				when "00101110111101" => data <= "111111";
				when "00101110111110" => data <= "100010";
				when "00101110111111" => data <= "111111";
				when "00101111000001" => data <= "111111";
				when "00101111000010" => data <= "100010";
				when "00101111000011" => data <= "111111";
				when "00110000001101" => data <= "111111";
				when "00110000001110" => data <= "110010";
				when "00110000001111" => data <= "111111";
				when "00110000010001" => data <= "111111";
				when "00110000010010" => data <= "110010";
				when "00110000010011" => data <= "111111";
				when "00110000010101" => data <= "111111";
				when "00110000010110" => data <= "110010";
				when "00110000010111" => data <= "111111";
				when "00110000011001" => data <= "111111";
				when "00110000011010" => data <= "110010";
				when "00110000011011" => data <= "111111";
				when "00110000011111" => data <= "111111";
				when "00110000100000" => data <= "110010";
				when "00110000100001" => data <= "111111";
				when "00110000100111" => data <= "111111";
				when "00110000101000" => data <= "110010";
				when "00110000101001" => data <= "111111";
				when "00110000101101" => data <= "111111";
				when "00110000101110" => data <= "110010";
				when "00110000101111" => data <= "111111";
				when "00110000110001" => data <= "111111";
				when "00110000110010" => data <= "110010";
				when "00110000110011" => data <= "111111";
				when "00110000110111" => data <= "111111";
				when "00110000111000" => data <= "110010";
				when "00110000111001" => data <= "111111";
				when "00110000111101" => data <= "111111";
				when "00110000111110" => data <= "110010";
				when "00110000111111" => data <= "111111";
				when "00110001000001" => data <= "111111";
				when "00110001000010" => data <= "110010";
				when "00110001000011" => data <= "111111";
				when "00110010001101" => data <= "111111";
				when "00110010001110" => data <= "110010";
				when "00110010001111" => data <= "111111";
				when "00110010010001" => data <= "111111";
				when "00110010010010" => data <= "110010";
				when "00110010010011" => data <= "111111";
				when "00110010010101" => data <= "111111";
				when "00110010010110" => data <= "110010";
				when "00110010010111" => data <= "111111";
				when "00110010011001" => data <= "111111";
				when "00110010011010" => data <= "110010";
				when "00110010011011" => data <= "111111";
				when "00110010011111" => data <= "111111";
				when "00110010100000" => data <= "110010";
				when "00110010100001" => data <= "111111";
				when "00110010100111" => data <= "111111";
				when "00110010101000" => data <= "110010";
				when "00110010101001" => data <= "111111";
				when "00110010101101" => data <= "111111";
				when "00110010101110" => data <= "110010";
				when "00110010101111" => data <= "111111";
				when "00110010110001" => data <= "111111";
				when "00110010110010" => data <= "110010";
				when "00110010110011" => data <= "111111";
				when "00110010110111" => data <= "111111";
				when "00110010111000" => data <= "110010";
				when "00110010111001" => data <= "111111";
				when "00110010111101" => data <= "111111";
				when "00110010111110" => data <= "110010";
				when "00110010111111" => data <= "111111";
				when "00110011000001" => data <= "111111";
				when "00110011000010" => data <= "110010";
				when "00110011000011" => data <= "111111";
				when "00110100001110" => data <= "111111";
				when "00110100010010" => data <= "111111";
				when "00110100010110" => data <= "111111";
				when "00110100011010" => data <= "111111";
				when "00110100100000" => data <= "111111";
				when "00110100101000" => data <= "111111";
				when "00110100101110" => data <= "111111";
				when "00110100110010" => data <= "111111";
				when "00110100111000" => data <= "111111";
				when "00110100111110" => data <= "111111";
				when "00110101000010" => data <= "111111";
				when "00111100011111" => data <= "010011";
				when "00111100100000" => data <= "010011";
				when "00111100110011" => data <= "010011";
				when "00111110011111" => data <= "010011";
				when "00111110100001" => data <= "010011";
				when "00111110100111" => data <= "010011";
				when "00111110101000" => data <= "010011";
				when "00111110101001" => data <= "010011";
				when "00111110101010" => data <= "010011";
				when "00111110101011" => data <= "010011";
				when "00111110110011" => data <= "010011";
				when "01000000011111" => data <= "010011";
				when "01000000100001" => data <= "010011";
				when "01000000100010" => data <= "010011";
				when "01000000100111" => data <= "010011";
				when "01000000101011" => data <= "010011";
				when "01000000110011" => data <= "010011";
				when "01000010011111" => data <= "010011";
				when "01000010100111" => data <= "010011";
				when "01000010101011" => data <= "010011";
				when "01000010110011" => data <= "010011";
				when "01000100011111" => data <= "010011";
				when "01000100100111" => data <= "010011";
				when "01000100101011" => data <= "010011";
				when "01000100110011" => data <= "010011";
				when "01000110011101" => data <= "010011";
				when "01000110011110" => data <= "010011";
				when "01000110011111" => data <= "010011";
				when "01000110100101" => data <= "010011";
				when "01000110100110" => data <= "010011";
				when "01000110100111" => data <= "010011";
				when "01000110101010" => data <= "010011";
				when "01000110101011" => data <= "010011";
				when "01000110110001" => data <= "010011";
				when "01000110110010" => data <= "010011";
				when "01000110110011" => data <= "010011";
				when "01001000011100" => data <= "110010";
				when "01001000011101" => data <= "111111";
				when "01001000011110" => data <= "010011";
				when "01001000011111" => data <= "110010";
				when "01001000100100" => data <= "010011";
				when "01001000100101" => data <= "111111";
				when "01001000100110" => data <= "010011";
				when "01001000100111" => data <= "010011";
				when "01001000101001" => data <= "111111";
				when "01001000101010" => data <= "010011";
				when "01001000101011" => data <= "010011";
				when "01001000110000" => data <= "110010";
				when "01001000110001" => data <= "111111";
				when "01001000110010" => data <= "010011";
				when "01001000110011" => data <= "110010";
				when "01001010011100" => data <= "100010";
				when "01001010011101" => data <= "110010";
				when "01001010011110" => data <= "110010";
				when "01001010011111" => data <= "100010";
				when "01001010100100" => data <= "100010";
				when "01001010100101" => data <= "110010";
				when "01001010100110" => data <= "110010";
				when "01001010100111" => data <= "100010";
				when "01001010101001" => data <= "100010";
				when "01001010101010" => data <= "110010";
				when "01001010101011" => data <= "100010";
				when "01001010110000" => data <= "100010";
				when "01001010110001" => data <= "110010";
				when "01001010110010" => data <= "110010";
				when "01001010110011" => data <= "100010";
				when "01001100011101" => data <= "100010";
				when "01001100011110" => data <= "100010";
				when "01001100100101" => data <= "100010";
				when "01001100100110" => data <= "100010";
				when "01001100101010" => data <= "100010";
				when "01001100110001" => data <= "100010";
				when "01001100110010" => data <= "100010";
				when "01011010001111" => data <= "111111";
				when "01011010010000" => data <= "111111";
				when "01011010010001" => data <= "111111";
				when "01011010010100" => data <= "111111";
				when "01011010010101" => data <= "111111";
				when "01011010010110" => data <= "111111";
				when "01011010011001" => data <= "111111";
				when "01011010011010" => data <= "111111";
				when "01011010011011" => data <= "111111";
				when "01011010011101" => data <= "111111";
				when "01011010011110" => data <= "111111";
				when "01011010011111" => data <= "111111";
				when "01011010100000" => data <= "111111";
				when "01011010100010" => data <= "111111";
				when "01011010100011" => data <= "111111";
				when "01011010100100" => data <= "111111";
				when "01011010100101" => data <= "111111";
				when "01011010101011" => data <= "111111";
				when "01011010101100" => data <= "111111";
				when "01011010101101" => data <= "111111";
				when "01011010101110" => data <= "111111";
				when "01011010110000" => data <= "111111";
				when "01011010110001" => data <= "111111";
				when "01011010110010" => data <= "111111";
				when "01011010110101" => data <= "111111";
				when "01011010110110" => data <= "111111";
				when "01011010111010" => data <= "111111";
				when "01011010111011" => data <= "111111";
				when "01011010111100" => data <= "111111";
				when "01011010111111" => data <= "111111";
				when "01011011000000" => data <= "111111";
				when "01011011000001" => data <= "111111";
				when "01011100001111" => data <= "111111";
				when "01011100010010" => data <= "111111";
				when "01011100010100" => data <= "111111";
				when "01011100010111" => data <= "111111";
				when "01011100011001" => data <= "111111";
				when "01011100011101" => data <= "111111";
				when "01011100100010" => data <= "111111";
				when "01011100101011" => data <= "111111";
				when "01011100110001" => data <= "111111";
				when "01011100110100" => data <= "111111";
				when "01011100110111" => data <= "111111";
				when "01011100111010" => data <= "111111";
				when "01011100111101" => data <= "111111";
				when "01011101000000" => data <= "111111";
				when "01011110001111" => data <= "111111";
				when "01011110010010" => data <= "111111";
				when "01011110010100" => data <= "111111";
				when "01011110010111" => data <= "111111";
				when "01011110011001" => data <= "111111";
				when "01011110011010" => data <= "111111";
				when "01011110011101" => data <= "111111";
				when "01011110011110" => data <= "111111";
				when "01011110011111" => data <= "111111";
				when "01011110100000" => data <= "111111";
				when "01011110100010" => data <= "111111";
				when "01011110100011" => data <= "111111";
				when "01011110100100" => data <= "111111";
				when "01011110100101" => data <= "111111";
				when "01011110101011" => data <= "111111";
				when "01011110101100" => data <= "111111";
				when "01011110101101" => data <= "111111";
				when "01011110101110" => data <= "111111";
				when "01011110110001" => data <= "111111";
				when "01011110110100" => data <= "111111";
				when "01011110110111" => data <= "111111";
				when "01011110111010" => data <= "111111";
				when "01011110111101" => data <= "111111";
				when "01011111000000" => data <= "111111";
				when "01100000001111" => data <= "111111";
				when "01100000010000" => data <= "111111";
				when "01100000010001" => data <= "111111";
				when "01100000010100" => data <= "111111";
				when "01100000010101" => data <= "111111";
				when "01100000010110" => data <= "111111";
				when "01100000011001" => data <= "111111";
				when "01100000100000" => data <= "111111";
				when "01100000100101" => data <= "111111";
				when "01100000101110" => data <= "111111";
				when "01100000110001" => data <= "111111";
				when "01100000110100" => data <= "111111";
				when "01100000110101" => data <= "111111";
				when "01100000110110" => data <= "111111";
				when "01100000110111" => data <= "111111";
				when "01100000111010" => data <= "111111";
				when "01100000111011" => data <= "111111";
				when "01100000111100" => data <= "111111";
				when "01100001000000" => data <= "111111";
				when "01100010001111" => data <= "111111";
				when "01100010010100" => data <= "111111";
				when "01100010010111" => data <= "111111";
				when "01100010011001" => data <= "111111";
				when "01100010100000" => data <= "111111";
				when "01100010100101" => data <= "111111";
				when "01100010101110" => data <= "111111";
				when "01100010110001" => data <= "111111";
				when "01100010110100" => data <= "111111";
				when "01100010110111" => data <= "111111";
				when "01100010111010" => data <= "111111";
				when "01100010111101" => data <= "111111";
				when "01100011000000" => data <= "111111";
				when "01100100001111" => data <= "111111";
				when "01100100010100" => data <= "111111";
				when "01100100010111" => data <= "111111";
				when "01100100011001" => data <= "111111";
				when "01100100011010" => data <= "111111";
				when "01100100011011" => data <= "111111";
				when "01100100011101" => data <= "111111";
				when "01100100011110" => data <= "111111";
				when "01100100011111" => data <= "111111";
				when "01100100100000" => data <= "111111";
				when "01100100100010" => data <= "111111";
				when "01100100100011" => data <= "111111";
				when "01100100100100" => data <= "111111";
				when "01100100100101" => data <= "111111";
				when "01100100101011" => data <= "111111";
				when "01100100101100" => data <= "111111";
				when "01100100101101" => data <= "111111";
				when "01100100101110" => data <= "111111";
				when "01100100110001" => data <= "111111";
				when "01100100110100" => data <= "111111";
				when "01100100110111" => data <= "111111";
				when "01100100111010" => data <= "111111";
				when "01100100111101" => data <= "111111";
				when "01100101000000" => data <= "111111";
				when others => data <= "000001";
			end case;
		end if; 
	end process; 
end;
