library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity alldig_disp is 
 	port(
		outglobal_o : in std_logic;
        digit : in std_logic_vector(3 downto 0);
		addr_x : in std_logic_vector(2 downto 0);
		addr_y : in std_logic_vector(2 downto 0);
		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
	);
end;

architecture sim of alldig_disp is
signal addr : std_logic_vector(9 downto 0);

begin
    addr (9 downto 6) <= digit;
	addr (5 downto 3) <= addr_x;
	addr (2 downto 0) <= addr_y;
	process(outglobal_o) begin
		if rising_edge(outglobal_o) then
			case addr is
                when "0000000000" => data <= "111111";
				when "0000000001" => data <= "111111";
				when "0000000010" => data <= "111111";
				when "0000000011" => data <= "111111";
				when "0000001000" => data <= "111111";
				when "0000001011" => data <= "111111";
				when "0000010000" => data <= "111111";
				when "0000010011" => data <= "111111";
				when "0000011000" => data <= "111111";
				when "0000011011" => data <= "111111";
				when "0000100000" => data <= "111111";
				when "0000100011" => data <= "111111";
				when "0000101000" => data <= "111111";
				when "0000101011" => data <= "111111";
				when "0000110000" => data <= "111111";
				when "0000110011" => data <= "111111";
				when "0000111000" => data <= "111111";
				when "0000111001" => data <= "111111";
				when "0000111010" => data <= "111111";
				when "0000111011" => data <= "111111";

                when "0001000010" => data <= "111111";
				when "0001001001" => data <= "111111";
				when "0001001010" => data <= "111111";
				when "0001010000" => data <= "111111";
				when "0001010010" => data <= "111111";
				when "0001011010" => data <= "111111";
				when "0001100010" => data <= "111111";
				when "0001101010" => data <= "111111";
				when "0001110010" => data <= "111111";
				when "0001111000" => data <= "111111";
				when "0001111001" => data <= "111111";
				when "0001111010" => data <= "111111";
				when "0001111011" => data <= "111111";

                when "0010000000" => data <= "111111";
				when "0010000001" => data <= "111111";
				when "0010000010" => data <= "111111";
				when "0010000011" => data <= "111111";
				when "0010001011" => data <= "111111";
				when "0010010011" => data <= "111111";
				when "0010011000" => data <= "111111";
				when "0010011001" => data <= "111111";
				when "0010011010" => data <= "111111";
				when "0010011011" => data <= "111111";
				when "0010100000" => data <= "111111";
				when "0010101000" => data <= "111111";
				when "0010110000" => data <= "111111";
				when "0010111000" => data <= "111111";
				when "0010111001" => data <= "111111";
				when "0010111010" => data <= "111111";
				when "0010111011" => data <= "111111";

                when "0011000000" => data <= "111111";
				when "0011000001" => data <= "111111";
				when "0011000010" => data <= "111111";
				when "0011000011" => data <= "111111";
				when "0011001011" => data <= "111111";
				when "0011010011" => data <= "111111";
				when "0011011001" => data <= "111111";
				when "0011011010" => data <= "111111";
				when "0011011011" => data <= "111111";
				when "0011100011" => data <= "111111";
				when "0011101011" => data <= "111111";
				when "0011110011" => data <= "111111";
				when "0011111000" => data <= "111111";
				when "0011111001" => data <= "111111";
				when "0011111010" => data <= "111111";
				when "0011111011" => data <= "111111";

                when "0100000000" => data <= "111111";
				when "0100000011" => data <= "111111";
				when "0100001000" => data <= "111111";
				when "0100001011" => data <= "111111";
				when "0100010000" => data <= "111111";
				when "0100010011" => data <= "111111";
				when "0100011000" => data <= "111111";
				when "0100011001" => data <= "111111";
				when "0100011010" => data <= "111111";
				when "0100011011" => data <= "111111";
				when "0100100011" => data <= "111111";
				when "0100101011" => data <= "111111";
				when "0100110011" => data <= "111111";
				when "0100111011" => data <= "111111";

                when "0101000000" => data <= "111111";
				when "0101000001" => data <= "111111";
				when "0101000010" => data <= "111111";
				when "0101000011" => data <= "111111";
				when "0101001000" => data <= "111111";
				when "0101010000" => data <= "111111";
				when "0101011000" => data <= "111111";
				when "0101011001" => data <= "111111";
				when "0101011010" => data <= "111111";
				when "0101011011" => data <= "111111";
				when "0101100011" => data <= "111111";
				when "0101101011" => data <= "111111";
				when "0101110011" => data <= "111111";
				when "0101111000" => data <= "111111";
				when "0101111001" => data <= "111111";
				when "0101111010" => data <= "111111";
				when "0101111011" => data <= "111111";

                when "0110000000" => data <= "111111";
				when "0110000001" => data <= "111111";
				when "0110000010" => data <= "111111";
				when "0110000011" => data <= "111111";
				when "0110001000" => data <= "111111";
				when "0110001011" => data <= "111111";
				when "0110010000" => data <= "111111";
				when "0110011000" => data <= "111111";
				when "0110011001" => data <= "111111";
				when "0110011010" => data <= "111111";
				when "0110011011" => data <= "111111";
				when "0110100000" => data <= "111111";
				when "0110100011" => data <= "111111";
				when "0110101000" => data <= "111111";
				when "0110101011" => data <= "111111";
				when "0110110000" => data <= "111111";
				when "0110110011" => data <= "111111";
				when "0110111000" => data <= "111111";
				when "0110111001" => data <= "111111";
				when "0110111010" => data <= "111111";
				when "0110111011" => data <= "111111";

                when "0111000000" => data <= "111111";
				when "0111000001" => data <= "111111";
				when "0111000010" => data <= "111111";
				when "0111000011" => data <= "111111";
				when "0111001011" => data <= "111111";
				when "0111010011" => data <= "111111";
				when "0111011011" => data <= "111111";
				when "0111100011" => data <= "111111";
				when "0111101011" => data <= "111111";
				when "0111110011" => data <= "111111";
				when "0111111011" => data <= "111111";

                when "1000000000" => data <= "111111";
				when "1000000001" => data <= "111111";
				when "1000000010" => data <= "111111";
				when "1000000011" => data <= "111111";
				when "1000001000" => data <= "111111";
				when "1000001011" => data <= "111111";
				when "1000010000" => data <= "111111";
				when "1000010011" => data <= "111111";
				when "1000011000" => data <= "111111";
				when "1000011001" => data <= "111111";
				when "1000011010" => data <= "111111";
				when "1000011011" => data <= "111111";
				when "1000100000" => data <= "111111";
				when "1000100011" => data <= "111111";
				when "1000101000" => data <= "111111";
				when "1000101011" => data <= "111111";
				when "1000110000" => data <= "111111";
				when "1000110011" => data <= "111111";
				when "1000111000" => data <= "111111";
				when "1000111001" => data <= "111111";
				when "1000111010" => data <= "111111";
				when "1000111011" => data <= "111111";

				when "1001000000" => data <= "111111";
				when "1001000001" => data <= "111111";
				when "1001000010" => data <= "111111";
				when "1001000011" => data <= "111111";
				when "1001001000" => data <= "111111";
				when "1001001011" => data <= "111111";
				when "1001010000" => data <= "111111";
				when "1001010011" => data <= "111111";
				when "1001011000" => data <= "111111";
				when "1001011001" => data <= "111111";
				when "1001011010" => data <= "111111";
				when "1001011011" => data <= "111111";
				when "1001100011" => data <= "111111";
				when "1001101011" => data <= "111111";
				when "1001110000" => data <= "111111";
				when "1001110011" => data <= "111111";
				when "1001111000" => data <= "111111";
				when "1001111001" => data <= "111111";
				when "1001111010" => data <= "111111";
				when "1001111011" => data <= "111111";
				when others => data <= "000001";
			end case;
		end if; 
	end process; 
end;