library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity rom is
                	port(
                		clk : in std_logic;
                		addr_x : in std_logic_vector(9 downto 0);
                		addr_y : in std_logic_vector(9 downto 0);
                		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
                	);
                end;

                architecture sim of rom is
                signal addr : std_logic_vector(18 downto 0);

                begin
                	addr (18 downto 10) <= addr_x;
                	addr (9 downto 0) <= addr_y;
                	process(clk) begin
                		if rising_edge(clk) then
                			case addr is
				when "000000000000000000" => data <= "010101";
				when "000000000000000001" => data <= "010101";
				when "000000000000000010" => data <= "010101";
				when "000000000000000011" => data <= "010101";
				when "000000000000000100" => data <= "010101";
				when "000000000000000101" => data <= "010101";
				when "000000000000000110" => data <= "010101";
				when "000000000000000111" => data <= "010101";
				when "000000000000001000" => data <= "010101";
				when "000000000000001001" => data <= "010101";
				when "000000000000001010" => data <= "010101";
				when "000000000000001011" => data <= "010101";
				when "000000000000001100" => data <= "010101";
				when "000000000000001101" => data <= "010101";
				when "000000000000001110" => data <= "010101";
				when "000000000000001111" => data <= "010101";
				when "000000000000010000" => data <= "010101";
				when "000000000000010001" => data <= "010101";
				when "000000000000010010" => data <= "010101";
				when "000000000000010011" => data <= "010101";
				when "000000000000010100" => data <= "010101";
				when "000000000000010101" => data <= "010101";
				when "000000000000010110" => data <= "010101";
				when "000000000000010111" => data <= "010101";
				when "000000000000011000" => data <= "010101";
				when "000000000000011001" => data <= "010101";
				when "000000000000011010" => data <= "010101";
				when "000000000000011011" => data <= "010101";
				when "000000000000011100" => data <= "010101";
				when "000000000000011101" => data <= "010101";
				when "000000000000011110" => data <= "010101";
				when "000000000000011111" => data <= "010101";
				when "000000000000100000" => data <= "010101";
				when "000000000000100001" => data <= "010101";
				when "000000000000100010" => data <= "010101";
				when "000000000000100011" => data <= "010101";
				when "000000000000100100" => data <= "010101";
				when "000000000000100101" => data <= "010101";
				when "000000000000100110" => data <= "010101";
				when "000000000000100111" => data <= "010101";
				when "000000000000101000" => data <= "010101";
				when "000000000000101001" => data <= "010101";
				when "000000000000101010" => data <= "010101";
				when "000000000000101011" => data <= "010101";
				when "000000000000101100" => data <= "010101";
				when "000000000000101101" => data <= "010101";
				when "000000000000101110" => data <= "010101";
				when "000000000000101111" => data <= "010101";
				when "000000000000110000" => data <= "010101";
				when "000000000000110001" => data <= "010101";
				when "000000000000110010" => data <= "010101";
				when "000000000000110011" => data <= "010101";
				when "000000000000110100" => data <= "010101";
				when "000000000000110101" => data <= "010101";
				when "000000000000110110" => data <= "010101";
				when "000000000000110111" => data <= "010101";
				when "000000000000111000" => data <= "010101";
				when "000000000000111001" => data <= "010101";
				when "000000000000111010" => data <= "010101";
				when "000000000000111011" => data <= "010101";
				when "000000000000111100" => data <= "010101";
				when "000000000000111101" => data <= "010101";
				when "000000000000111110" => data <= "010101";
				when "000000000000111111" => data <= "010101";
				when "000000000001000000" => data <= "010101";
				when "000000000001000001" => data <= "010101";
				when "000000000001000010" => data <= "010101";
				when "000000000001000011" => data <= "010101";
				when "000000000001000100" => data <= "010101";
				when "000000000001000101" => data <= "010101";
				when "000000000001000110" => data <= "010101";
				when "000000000001000111" => data <= "010101";
				when "000000000001001000" => data <= "010101";
				when "000000000001001001" => data <= "010101";
				when "000000000001001010" => data <= "010101";
				when "000000000001001011" => data <= "010101";
				when "000000000001001100" => data <= "010101";
				when "000000000001001101" => data <= "010101";
				when "000000000001001110" => data <= "010101";
				when "000000000001001111" => data <= "010101";
				when "000000000001010000" => data <= "010101";
				when "000000000001010001" => data <= "010101";
				when "000000000001010010" => data <= "010101";
				when "000000000001010011" => data <= "010101";
				when "000000000001010100" => data <= "010101";
				when "000000000001010101" => data <= "010101";
				when "000000000001010110" => data <= "010101";
				when "000000000001010111" => data <= "010101";
				when "000000000001011000" => data <= "010101";
				when "000000000001011001" => data <= "010101";
				when "000000000001011010" => data <= "010101";
				when "000000000001011011" => data <= "010101";
				when "000000000001011100" => data <= "010101";
				when "000000000001011101" => data <= "010101";
				when "000000000001011110" => data <= "010101";
				when "000000000001011111" => data <= "010101";
				when "000000000001100000" => data <= "010101";
				when "000000000001100001" => data <= "010101";
				when "000000000001100010" => data <= "010101";
				when "000000000001100011" => data <= "010101";
				when "000000000001100100" => data <= "010101";
				when "000000000001100101" => data <= "010101";
				when "000000000001100110" => data <= "010101";
				when "000000000001100111" => data <= "010101";
				when "000000000001101000" => data <= "010101";
				when "000000000001101001" => data <= "010101";
				when "000000000001101010" => data <= "010101";
				when "000000000001101011" => data <= "010101";
				when "000000000001101100" => data <= "010101";
				when "000000000001101101" => data <= "010101";
				when "000000000001101110" => data <= "010101";
				when "000000000001101111" => data <= "010101";
				when "000000000001110000" => data <= "010101";
				when "000000000001110001" => data <= "010101";
				when "000000000001110010" => data <= "010101";
				when "000000000001110011" => data <= "010101";
				when "000000000001110100" => data <= "010101";
				when "000000000001110101" => data <= "010101";
				when "000000000001110110" => data <= "010101";
				when "000000000001110111" => data <= "010101";
				when "000000000001111000" => data <= "010101";
				when "000000000001111001" => data <= "010101";
				when "000000000001111010" => data <= "010101";
				when "000000000001111011" => data <= "010101";
				when "000000000001111100" => data <= "010101";
				when "000000000001111101" => data <= "010101";
				when "000000000001111110" => data <= "010101";
				when "000000000001111111" => data <= "010101";
				when "000000000010000000" => data <= "010101";
				when "000000000010000001" => data <= "010101";
				when "000000000010000010" => data <= "010101";
				when "000000000010000011" => data <= "010101";
				when "000000000010000100" => data <= "010101";
				when "000000000010000101" => data <= "010101";
				when "000000000010000110" => data <= "010101";
				when "000000000010000111" => data <= "010101";
				when "000000000010001000" => data <= "010101";
				when "000000000010001001" => data <= "010101";
				when "000000000010001010" => data <= "010101";
				when "000000000010001011" => data <= "010101";
				when "000000000010001100" => data <= "010101";
				when "000000000010001101" => data <= "010101";
				when "000000000010001110" => data <= "010101";
				when "000000000010001111" => data <= "010101";
				when "000000000010010000" => data <= "010101";
				when "000000000010010001" => data <= "010101";
				when "000000000010010010" => data <= "010101";
				when "000000000010010011" => data <= "010101";
				when "000000000010010100" => data <= "010101";
				when "000000000010010101" => data <= "010101";
				when "000000000010010110" => data <= "010101";
				when "000000000010010111" => data <= "010101";
				when "000000000010011000" => data <= "010101";
				when "000000000010011001" => data <= "010101";
				when "000000000010011010" => data <= "010101";
				when "000000000010011011" => data <= "010101";
				when "000000000010011100" => data <= "010101";
				when "000000000010011101" => data <= "010101";
				when "000000000010011110" => data <= "010101";
				when "000000000010011111" => data <= "010101";
				when "000000001000000000" => data <= "010101";
				when "000000001000000001" => data <= "010101";
				when "000000001000000010" => data <= "010101";
				when "000000001000000011" => data <= "010101";
				when "000000001000000100" => data <= "010101";
				when "000000001000000101" => data <= "010101";
				when "000000001000000110" => data <= "010101";
				when "000000001000000111" => data <= "010101";
				when "000000001000001000" => data <= "010101";
				when "000000001000001001" => data <= "010101";
				when "000000001000001010" => data <= "010101";
				when "000000001000001011" => data <= "010101";
				when "000000001000001100" => data <= "010101";
				when "000000001000001101" => data <= "010101";
				when "000000001000001110" => data <= "010101";
				when "000000001000001111" => data <= "010101";
				when "000000001000010000" => data <= "010101";
				when "000000001000010001" => data <= "010101";
				when "000000001000010010" => data <= "010101";
				when "000000001000010011" => data <= "010101";
				when "000000001000010100" => data <= "010101";
				when "000000001000010101" => data <= "010101";
				when "000000001000010110" => data <= "010101";
				when "000000001000010111" => data <= "010101";
				when "000000001000011000" => data <= "010101";
				when "000000001000011001" => data <= "010101";
				when "000000001000011010" => data <= "010101";
				when "000000001000011011" => data <= "010101";
				when "000000001000011100" => data <= "010101";
				when "000000001000011101" => data <= "010101";
				when "000000001000011110" => data <= "010101";
				when "000000001000011111" => data <= "010101";
				when "000000001000100000" => data <= "010101";
				when "000000001000100001" => data <= "010101";
				when "000000001000100010" => data <= "010101";
				when "000000001000100011" => data <= "010101";
				when "000000001000100100" => data <= "010101";
				when "000000001000100101" => data <= "010101";
				when "000000001000100110" => data <= "010101";
				when "000000001000100111" => data <= "010101";
				when "000000001000101000" => data <= "010101";
				when "000000001000101001" => data <= "010101";
				when "000000001000101010" => data <= "010101";
				when "000000001000101011" => data <= "010101";
				when "000000001000101100" => data <= "010101";
				when "000000001000101101" => data <= "010101";
				when "000000001000101110" => data <= "010101";
				when "000000001000101111" => data <= "010101";
				when "000000001000110000" => data <= "010101";
				when "000000001000110001" => data <= "010101";
				when "000000001000110010" => data <= "010101";
				when "000000001000110011" => data <= "010101";
				when "000000001000110100" => data <= "010101";
				when "000000001000110101" => data <= "010101";
				when "000000001000110110" => data <= "010101";
				when "000000001000110111" => data <= "010101";
				when "000000001000111000" => data <= "010101";
				when "000000001000111001" => data <= "010101";
				when "000000001000111010" => data <= "010101";
				when "000000001000111011" => data <= "010101";
				when "000000001000111100" => data <= "010101";
				when "000000001000111101" => data <= "010101";
				when "000000001000111110" => data <= "010101";
				when "000000001000111111" => data <= "010101";
				when "000000001001000000" => data <= "010101";
				when "000000001001000001" => data <= "010101";
				when "000000001001000010" => data <= "010101";
				when "000000001001000011" => data <= "010101";
				when "000000001001000100" => data <= "010101";
				when "000000001001000101" => data <= "010101";
				when "000000001001000110" => data <= "010101";
				when "000000001001000111" => data <= "010101";
				when "000000001001001000" => data <= "010101";
				when "000000001001001001" => data <= "010101";
				when "000000001001001010" => data <= "010101";
				when "000000001001001011" => data <= "010101";
				when "000000001001001100" => data <= "010101";
				when "000000001001001101" => data <= "010101";
				when "000000001001001110" => data <= "010101";
				when "000000001001001111" => data <= "010101";
				when "000000001001010000" => data <= "010101";
				when "000000001001010001" => data <= "010101";
				when "000000001001010010" => data <= "010101";
				when "000000001001010011" => data <= "010101";
				when "000000001001010100" => data <= "010101";
				when "000000001001010101" => data <= "010101";
				when "000000001001010110" => data <= "010101";
				when "000000001001010111" => data <= "010101";
				when "000000001001011000" => data <= "010101";
				when "000000001001011001" => data <= "010101";
				when "000000001001011010" => data <= "010101";
				when "000000001001011011" => data <= "010101";
				when "000000001001011100" => data <= "010101";
				when "000000001001011101" => data <= "010101";
				when "000000001001011110" => data <= "010101";
				when "000000001001011111" => data <= "010101";
				when "000000001001100000" => data <= "010101";
				when "000000001001100001" => data <= "010101";
				when "000000001001100010" => data <= "010101";
				when "000000001001100011" => data <= "010101";
				when "000000001001100100" => data <= "010101";
				when "000000001001100101" => data <= "010101";
				when "000000001001100110" => data <= "010101";
				when "000000001001100111" => data <= "010101";
				when "000000001001101000" => data <= "010101";
				when "000000001001101001" => data <= "010101";
				when "000000001001101010" => data <= "010101";
				when "000000001001101011" => data <= "010101";
				when "000000001001101100" => data <= "010101";
				when "000000001001101101" => data <= "010101";
				when "000000001001101110" => data <= "010101";
				when "000000001001101111" => data <= "010101";
				when "000000001001110000" => data <= "010101";
				when "000000001001110001" => data <= "010101";
				when "000000001001110010" => data <= "010101";
				when "000000001001110011" => data <= "010101";
				when "000000001001110100" => data <= "010101";
				when "000000001001110101" => data <= "010101";
				when "000000001001110110" => data <= "010101";
				when "000000001001110111" => data <= "010101";
				when "000000001001111000" => data <= "010101";
				when "000000001001111001" => data <= "010101";
				when "000000001001111010" => data <= "010101";
				when "000000001001111011" => data <= "010101";
				when "000000001001111100" => data <= "010101";
				when "000000001001111101" => data <= "010101";
				when "000000001001111110" => data <= "010101";
				when "000000001001111111" => data <= "010101";
				when "000000001010000000" => data <= "010101";
				when "000000001010000001" => data <= "010101";
				when "000000001010000010" => data <= "010101";
				when "000000001010000011" => data <= "010101";
				when "000000001010000100" => data <= "010101";
				when "000000001010000101" => data <= "010101";
				when "000000001010000110" => data <= "010101";
				when "000000001010000111" => data <= "010101";
				when "000000001010001000" => data <= "010101";
				when "000000001010001001" => data <= "010101";
				when "000000001010001010" => data <= "010101";
				when "000000001010001011" => data <= "010101";
				when "000000001010001100" => data <= "010101";
				when "000000001010001101" => data <= "010101";
				when "000000001010001110" => data <= "010101";
				when "000000001010001111" => data <= "010101";
				when "000000001010010000" => data <= "010101";
				when "000000001010010001" => data <= "010101";
				when "000000001010010010" => data <= "010101";
				when "000000001010010011" => data <= "010101";
				when "000000001010010100" => data <= "010101";
				when "000000001010010101" => data <= "010101";
				when "000000001010010110" => data <= "010101";
				when "000000001010010111" => data <= "010101";
				when "000000001010011000" => data <= "010101";
				when "000000001010011001" => data <= "010101";
				when "000000001010011010" => data <= "010101";
				when "000000001010011011" => data <= "010101";
				when "000000001010011100" => data <= "010101";
				when "000000001010011101" => data <= "010101";
				when "000000001010011110" => data <= "010101";
				when "000000001010011111" => data <= "010101";
				when "000000010000000000" => data <= "010101";
				when "000000010000000001" => data <= "010101";
				when "000000010000000010" => data <= "010101";
				when "000000010000000011" => data <= "010101";
				when "000000010000000100" => data <= "010101";
				when "000000010000000101" => data <= "010101";
				when "000000010000000110" => data <= "010101";
				when "000000010000000111" => data <= "010101";
				when "000000010000001000" => data <= "010101";
				when "000000010000001001" => data <= "010101";
				when "000000010000001010" => data <= "010101";
				when "000000010000001011" => data <= "010101";
				when "000000010000001100" => data <= "010101";
				when "000000010000001101" => data <= "010101";
				when "000000010000001110" => data <= "010101";
				when "000000010000001111" => data <= "010101";
				when "000000010000010000" => data <= "010101";
				when "000000010000010001" => data <= "010101";
				when "000000010000010010" => data <= "010101";
				when "000000010000010011" => data <= "010101";
				when "000000010000010100" => data <= "010101";
				when "000000010000010101" => data <= "010101";
				when "000000010000010110" => data <= "010101";
				when "000000010000010111" => data <= "010101";
				when "000000010000011000" => data <= "010101";
				when "000000010000011001" => data <= "010101";
				when "000000010000011010" => data <= "010101";
				when "000000010000011011" => data <= "010101";
				when "000000010000011100" => data <= "010101";
				when "000000010000011101" => data <= "010101";
				when "000000010000011110" => data <= "010101";
				when "000000010000011111" => data <= "010101";
				when "000000010000100000" => data <= "010101";
				when "000000010000100001" => data <= "010101";
				when "000000010000100010" => data <= "010101";
				when "000000010000100011" => data <= "010101";
				when "000000010000100100" => data <= "010101";
				when "000000010000100101" => data <= "010101";
				when "000000010000100110" => data <= "010101";
				when "000000010000100111" => data <= "010101";
				when "000000010000101000" => data <= "010101";
				when "000000010000101001" => data <= "010101";
				when "000000010000101010" => data <= "010101";
				when "000000010000101011" => data <= "010101";
				when "000000010000101100" => data <= "010101";
				when "000000010000101101" => data <= "010101";
				when "000000010000101110" => data <= "010101";
				when "000000010000101111" => data <= "010101";
				when "000000010000110000" => data <= "010101";
				when "000000010000110001" => data <= "010101";
				when "000000010000110010" => data <= "010101";
				when "000000010000110011" => data <= "010101";
				when "000000010000110100" => data <= "010101";
				when "000000010000110101" => data <= "010101";
				when "000000010000110110" => data <= "010101";
				when "000000010000110111" => data <= "010101";
				when "000000010000111000" => data <= "010101";
				when "000000010000111001" => data <= "010101";
				when "000000010000111010" => data <= "010101";
				when "000000010000111011" => data <= "010101";
				when "000000010000111100" => data <= "010101";
				when "000000010000111101" => data <= "010101";
				when "000000010000111110" => data <= "010101";
				when "000000010000111111" => data <= "010101";
				when "000000010001000000" => data <= "010101";
				when "000000010001000001" => data <= "010101";
				when "000000010001000010" => data <= "010101";
				when "000000010001000011" => data <= "010101";
				when "000000010001000100" => data <= "010101";
				when "000000010001000101" => data <= "010101";
				when "000000010001000110" => data <= "010101";
				when "000000010001000111" => data <= "010101";
				when "000000010001001000" => data <= "010101";
				when "000000010001001001" => data <= "010101";
				when "000000010001001010" => data <= "010101";
				when "000000010001001011" => data <= "010101";
				when "000000010001001100" => data <= "010101";
				when "000000010001001101" => data <= "010101";
				when "000000010001001110" => data <= "010101";
				when "000000010001001111" => data <= "010101";
				when "000000010001010000" => data <= "010101";
				when "000000010001010001" => data <= "010101";
				when "000000010001010010" => data <= "010101";
				when "000000010001010011" => data <= "010101";
				when "000000010001010100" => data <= "010101";
				when "000000010001010101" => data <= "010101";
				when "000000010001010110" => data <= "010101";
				when "000000010001010111" => data <= "010101";
				when "000000010001011000" => data <= "010101";
				when "000000010001011001" => data <= "010101";
				when "000000010001011010" => data <= "010101";
				when "000000010001011011" => data <= "010101";
				when "000000010001011100" => data <= "010101";
				when "000000010001011101" => data <= "010101";
				when "000000010001011110" => data <= "010101";
				when "000000010001011111" => data <= "010101";
				when "000000010001100000" => data <= "010101";
				when "000000010001100001" => data <= "010101";
				when "000000010001100010" => data <= "010101";
				when "000000010001100011" => data <= "010101";
				when "000000010001100100" => data <= "010101";
				when "000000010001100101" => data <= "010101";
				when "000000010001100110" => data <= "010101";
				when "000000010001100111" => data <= "010101";
				when "000000010001101000" => data <= "010101";
				when "000000010001101001" => data <= "010101";
				when "000000010001101010" => data <= "010101";
				when "000000010001101011" => data <= "010101";
				when "000000010001101100" => data <= "010101";
				when "000000010001101101" => data <= "010101";
				when "000000010001101110" => data <= "010101";
				when "000000010001101111" => data <= "010101";
				when "000000010001110000" => data <= "010101";
				when "000000010001110001" => data <= "010101";
				when "000000010001110010" => data <= "010101";
				when "000000010001110011" => data <= "010101";
				when "000000010001110100" => data <= "010101";
				when "000000010001110101" => data <= "010101";
				when "000000010001110110" => data <= "010101";
				when "000000010001110111" => data <= "010101";
				when "000000010001111000" => data <= "010101";
				when "000000010001111001" => data <= "010101";
				when "000000010001111010" => data <= "010101";
				when "000000010001111011" => data <= "010101";
				when "000000010001111100" => data <= "010101";
				when "000000010001111101" => data <= "010101";
				when "000000010001111110" => data <= "010101";
				when "000000010001111111" => data <= "010101";
				when "000000010010000000" => data <= "010101";
				when "000000010010000001" => data <= "010101";
				when "000000010010000010" => data <= "010101";
				when "000000010010000011" => data <= "010101";
				when "000000010010000100" => data <= "010101";
				when "000000010010000101" => data <= "010101";
				when "000000010010000110" => data <= "010101";
				when "000000010010000111" => data <= "010101";
				when "000000010010001000" => data <= "010101";
				when "000000010010001001" => data <= "010101";
				when "000000010010001010" => data <= "010101";
				when "000000010010001011" => data <= "010101";
				when "000000010010001100" => data <= "010101";
				when "000000010010001101" => data <= "010101";
				when "000000010010001110" => data <= "010101";
				when "000000010010001111" => data <= "010101";
				when "000000010010010000" => data <= "010101";
				when "000000010010010001" => data <= "010101";
				when "000000010010010010" => data <= "010101";
				when "000000010010010011" => data <= "010101";
				when "000000010010010100" => data <= "010101";
				when "000000010010010101" => data <= "010101";
				when "000000010010010110" => data <= "010101";
				when "000000010010010111" => data <= "010101";
				when "000000010010011000" => data <= "010101";
				when "000000010010011001" => data <= "010101";
				when "000000010010011010" => data <= "010101";
				when "000000010010011011" => data <= "010101";
				when "000000010010011100" => data <= "010101";
				when "000000010010011101" => data <= "010101";
				when "000000010010011110" => data <= "010101";
				when "000000010010011111" => data <= "010101";
				when "000000011000000000" => data <= "010101";
				when "000000011000000001" => data <= "010101";
				when "000000011000000010" => data <= "010101";
				when "000000011000000011" => data <= "010101";
				when "000000011000000100" => data <= "010101";
				when "000000011000000101" => data <= "010101";
				when "000000011000000110" => data <= "010101";
				when "000000011000000111" => data <= "010101";
				when "000000011000001000" => data <= "010101";
				when "000000011000001001" => data <= "010101";
				when "000000011000001010" => data <= "010101";
				when "000000011000001011" => data <= "010101";
				when "000000011000001100" => data <= "010101";
				when "000000011000001101" => data <= "010101";
				when "000000011000001110" => data <= "010101";
				when "000000011000001111" => data <= "010101";
				when "000000011000010000" => data <= "010101";
				when "000000011000010001" => data <= "010101";
				when "000000011000010010" => data <= "010101";
				when "000000011000010011" => data <= "010101";
				when "000000011000010100" => data <= "010101";
				when "000000011000010101" => data <= "010101";
				when "000000011000010110" => data <= "010101";
				when "000000011000010111" => data <= "010101";
				when "000000011000011000" => data <= "010101";
				when "000000011000011001" => data <= "010101";
				when "000000011000011010" => data <= "010101";
				when "000000011000011011" => data <= "010101";
				when "000000011000011100" => data <= "010101";
				when "000000011000011101" => data <= "010101";
				when "000000011000011110" => data <= "010101";
				when "000000011000011111" => data <= "010101";
				when "000000011000100000" => data <= "010101";
				when "000000011000100001" => data <= "010101";
				when "000000011000100010" => data <= "010101";
				when "000000011000100011" => data <= "010101";
				when "000000011000100100" => data <= "010101";
				when "000000011000100101" => data <= "010101";
				when "000000011000100110" => data <= "010101";
				when "000000011000100111" => data <= "010101";
				when "000000011000101000" => data <= "010101";
				when "000000011000101001" => data <= "010101";
				when "000000011000101010" => data <= "010101";
				when "000000011000101011" => data <= "010101";
				when "000000011000101100" => data <= "010101";
				when "000000011000101101" => data <= "010101";
				when "000000011000101110" => data <= "010101";
				when "000000011000101111" => data <= "010101";
				when "000000011000110000" => data <= "010101";
				when "000000011000110001" => data <= "010101";
				when "000000011000110010" => data <= "010101";
				when "000000011000110011" => data <= "010101";
				when "000000011000110100" => data <= "010101";
				when "000000011000110101" => data <= "010101";
				when "000000011000110110" => data <= "010101";
				when "000000011000110111" => data <= "010101";
				when "000000011000111000" => data <= "010101";
				when "000000011000111001" => data <= "010101";
				when "000000011000111010" => data <= "010101";
				when "000000011000111011" => data <= "010101";
				when "000000011000111100" => data <= "010101";
				when "000000011000111101" => data <= "010101";
				when "000000011000111110" => data <= "010101";
				when "000000011000111111" => data <= "010101";
				when "000000011001000000" => data <= "010101";
				when "000000011001000001" => data <= "010101";
				when "000000011001000010" => data <= "010101";
				when "000000011001000011" => data <= "010101";
				when "000000011001000100" => data <= "010101";
				when "000000011001000101" => data <= "010101";
				when "000000011001000110" => data <= "010101";
				when "000000011001000111" => data <= "010101";
				when "000000011001001000" => data <= "010101";
				when "000000011001001001" => data <= "010101";
				when "000000011001001010" => data <= "010101";
				when "000000011001001011" => data <= "010101";
				when "000000011001001100" => data <= "010101";
				when "000000011001001101" => data <= "010101";
				when "000000011001001110" => data <= "010101";
				when "000000011001001111" => data <= "010101";
				when "000000011001010000" => data <= "010101";
				when "000000011001010001" => data <= "010101";
				when "000000011001010010" => data <= "010101";
				when "000000011001010011" => data <= "010101";
				when "000000011001010100" => data <= "010101";
				when "000000011001010101" => data <= "010101";
				when "000000011001010110" => data <= "010101";
				when "000000011001010111" => data <= "010101";
				when "000000011001011000" => data <= "010101";
				when "000000011001011001" => data <= "010101";
				when "000000011001011010" => data <= "010101";
				when "000000011001011011" => data <= "010101";
				when "000000011001011100" => data <= "010101";
				when "000000011001011101" => data <= "010101";
				when "000000011001011110" => data <= "010101";
				when "000000011001011111" => data <= "010101";
				when "000000011001100000" => data <= "010101";
				when "000000011001100001" => data <= "010101";
				when "000000011001100010" => data <= "010101";
				when "000000011001100011" => data <= "010101";
				when "000000011001100100" => data <= "010101";
				when "000000011001100101" => data <= "010101";
				when "000000011001100110" => data <= "010101";
				when "000000011001100111" => data <= "010101";
				when "000000011001101000" => data <= "010101";
				when "000000011001101001" => data <= "010101";
				when "000000011001101010" => data <= "010101";
				when "000000011001101011" => data <= "010101";
				when "000000011001101100" => data <= "010101";
				when "000000011001101101" => data <= "010101";
				when "000000011001101110" => data <= "010101";
				when "000000011001101111" => data <= "010101";
				when "000000011001110000" => data <= "010101";
				when "000000011001110001" => data <= "010101";
				when "000000011001110010" => data <= "010101";
				when "000000011001110011" => data <= "010101";
				when "000000011001110100" => data <= "010101";
				when "000000011001110101" => data <= "010101";
				when "000000011001110110" => data <= "010101";
				when "000000011001110111" => data <= "010101";
				when "000000011001111000" => data <= "010101";
				when "000000011001111001" => data <= "010101";
				when "000000011001111010" => data <= "010101";
				when "000000011001111011" => data <= "010101";
				when "000000011001111100" => data <= "010101";
				when "000000011001111101" => data <= "010101";
				when "000000011001111110" => data <= "010101";
				when "000000011001111111" => data <= "010101";
				when "000000011010000000" => data <= "010101";
				when "000000011010000001" => data <= "010101";
				when "000000011010000010" => data <= "010101";
				when "000000011010000011" => data <= "010101";
				when "000000011010000100" => data <= "010101";
				when "000000011010000101" => data <= "010101";
				when "000000011010000110" => data <= "010101";
				when "000000011010000111" => data <= "010101";
				when "000000011010001000" => data <= "010101";
				when "000000011010001001" => data <= "010101";
				when "000000011010001010" => data <= "010101";
				when "000000011010001011" => data <= "010101";
				when "000000011010001100" => data <= "010101";
				when "000000011010001101" => data <= "010101";
				when "000000011010001110" => data <= "010101";
				when "000000011010001111" => data <= "010101";
				when "000000011010010000" => data <= "010101";
				when "000000011010010001" => data <= "010101";
				when "000000011010010010" => data <= "010101";
				when "000000011010010011" => data <= "010101";
				when "000000011010010100" => data <= "010101";
				when "000000011010010101" => data <= "010101";
				when "000000011010010110" => data <= "010101";
				when "000000011010010111" => data <= "010101";
				when "000000011010011000" => data <= "010101";
				when "000000011010011001" => data <= "010101";
				when "000000011010011010" => data <= "010101";
				when "000000011010011011" => data <= "010101";
				when "000000011010011100" => data <= "010101";
				when "000000011010011101" => data <= "010101";
				when "000000011010011110" => data <= "010101";
				when "000000011010011111" => data <= "010101";
				when "000000100000000000" => data <= "000000";
				when "000000100000000001" => data <= "000000";
				when "000000100000000010" => data <= "000000";
				when "000000100000000011" => data <= "000000";
				when "000000100000000100" => data <= "000000";
				when "000000100000000101" => data <= "000000";
				when "000000100000000110" => data <= "000000";
				when "000000100000000111" => data <= "000000";
				when "000000100000001000" => data <= "000000";
				when "000000100000001001" => data <= "000000";
				when "000000100000001010" => data <= "000000";
				when "000000100000001011" => data <= "000000";
				when "000000100000001100" => data <= "000000";
				when "000000100000001101" => data <= "000000";
				when "000000100000001110" => data <= "000000";
				when "000000100000001111" => data <= "000000";
				when "000000100000010000" => data <= "000000";
				when "000000100000010001" => data <= "000000";
				when "000000100000010010" => data <= "000000";
				when "000000100000010011" => data <= "000000";
				when "000000100000010100" => data <= "000000";
				when "000000100000010101" => data <= "000000";
				when "000000100000010110" => data <= "000000";
				when "000000100000010111" => data <= "000000";
				when "000000100000011000" => data <= "000000";
				when "000000100000011001" => data <= "000000";
				when "000000100000011010" => data <= "000000";
				when "000000100000011011" => data <= "000000";
				when "000000100000011100" => data <= "000000";
				when "000000100000011101" => data <= "000000";
				when "000000100000011110" => data <= "000000";
				when "000000100000011111" => data <= "000000";
				when "000000100000100000" => data <= "000000";
				when "000000100000100001" => data <= "000000";
				when "000000100000100010" => data <= "000000";
				when "000000100000100011" => data <= "000000";
				when "000000100000100100" => data <= "000000";
				when "000000100000100101" => data <= "000000";
				when "000000100000100110" => data <= "000000";
				when "000000100000100111" => data <= "000000";
				when "000000100000101000" => data <= "000000";
				when "000000100000101001" => data <= "000000";
				when "000000100000101010" => data <= "000000";
				when "000000100000101011" => data <= "000000";
				when "000000100000101100" => data <= "000000";
				when "000000100000101101" => data <= "000000";
				when "000000100000101110" => data <= "000000";
				when "000000100000101111" => data <= "000000";
				when "000000100000110000" => data <= "000000";
				when "000000100000110001" => data <= "000000";
				when "000000100000110010" => data <= "000000";
				when "000000100000110011" => data <= "000000";
				when "000000100000110100" => data <= "000000";
				when "000000100000110101" => data <= "000000";
				when "000000100000110110" => data <= "000000";
				when "000000100000110111" => data <= "000000";
				when "000000100000111000" => data <= "000000";
				when "000000100000111001" => data <= "000000";
				when "000000100000111010" => data <= "000000";
				when "000000100000111011" => data <= "000000";
				when "000000100000111100" => data <= "000000";
				when "000000100000111101" => data <= "000000";
				when "000000100000111110" => data <= "000000";
				when "000000100000111111" => data <= "000000";
				when "000000100001000000" => data <= "000000";
				when "000000100001000001" => data <= "000000";
				when "000000100001000010" => data <= "000000";
				when "000000100001000011" => data <= "000000";
				when "000000100001000100" => data <= "000000";
				when "000000100001000101" => data <= "000000";
				when "000000100001000110" => data <= "000000";
				when "000000100001000111" => data <= "000000";
				when "000000100001001000" => data <= "000000";
				when "000000100001001001" => data <= "000000";
				when "000000100001001010" => data <= "000000";
				when "000000100001001011" => data <= "000000";
				when "000000100001001100" => data <= "000000";
				when "000000100001001101" => data <= "000000";
				when "000000100001001110" => data <= "000000";
				when "000000100001001111" => data <= "000000";
				when "000000100001010000" => data <= "000000";
				when "000000100001010001" => data <= "000000";
				when "000000100001010010" => data <= "000000";
				when "000000100001010011" => data <= "000000";
				when "000000100001010100" => data <= "000000";
				when "000000100001010101" => data <= "000000";
				when "000000100001010110" => data <= "000000";
				when "000000100001010111" => data <= "000000";
				when "000000100001011000" => data <= "000000";
				when "000000100001011001" => data <= "000000";
				when "000000100001011010" => data <= "000000";
				when "000000100001011011" => data <= "000000";
				when "000000100001011100" => data <= "000000";
				when "000000100001011101" => data <= "000000";
				when "000000100001011110" => data <= "000000";
				when "000000100001011111" => data <= "000000";
				when "000000100001100000" => data <= "000000";
				when "000000100001100001" => data <= "000000";
				when "000000100001100010" => data <= "000000";
				when "000000100001100011" => data <= "000000";
				when "000000100001100100" => data <= "000000";
				when "000000100001100101" => data <= "000000";
				when "000000100001100110" => data <= "000000";
				when "000000100001100111" => data <= "000000";
				when "000000100001101000" => data <= "000000";
				when "000000100001101001" => data <= "000000";
				when "000000100001101010" => data <= "000000";
				when "000000100001101011" => data <= "000000";
				when "000000100001101100" => data <= "000000";
				when "000000100001101101" => data <= "000000";
				when "000000100001101110" => data <= "000000";
				when "000000100001101111" => data <= "000000";
				when "000000100001110000" => data <= "000000";
				when "000000100001110001" => data <= "000000";
				when "000000100001110010" => data <= "000000";
				when "000000100001110011" => data <= "000000";
				when "000000100001110100" => data <= "000000";
				when "000000100001110101" => data <= "000000";
				when "000000100001110110" => data <= "000000";
				when "000000100001110111" => data <= "000000";
				when "000000100001111000" => data <= "000000";
				when "000000100001111001" => data <= "000000";
				when "000000100001111010" => data <= "000000";
				when "000000100001111011" => data <= "000000";
				when "000000100001111100" => data <= "000000";
				when "000000100001111101" => data <= "000000";
				when "000000100001111110" => data <= "000000";
				when "000000100001111111" => data <= "000000";
				when "000000100010000000" => data <= "000000";
				when "000000100010000001" => data <= "000000";
				when "000000100010000010" => data <= "000000";
				when "000000100010000011" => data <= "000000";
				when "000000100010000100" => data <= "000000";
				when "000000100010000101" => data <= "000000";
				when "000000100010000110" => data <= "000000";
				when "000000100010000111" => data <= "000000";
				when "000000100010001000" => data <= "000000";
				when "000000100010001001" => data <= "000000";
				when "000000100010001010" => data <= "000000";
				when "000000100010001011" => data <= "000000";
				when "000000100010001100" => data <= "000000";
				when "000000100010001101" => data <= "000000";
				when "000000100010001110" => data <= "000000";
				when "000000100010001111" => data <= "000000";
				when "000000100010010000" => data <= "000000";
				when "000000100010010001" => data <= "000000";
				when "000000100010010010" => data <= "000000";
				when "000000100010010011" => data <= "000000";
				when "000000100010010100" => data <= "000000";
				when "000000100010010101" => data <= "000000";
				when "000000100010010110" => data <= "000000";
				when "000000100010010111" => data <= "000000";
				when "000000100010011000" => data <= "000000";
				when "000000100010011001" => data <= "000000";
				when "000000100010011010" => data <= "000000";
				when "000000100010011011" => data <= "000000";
				when "000000100010011100" => data <= "000000";
				when "000000100010011101" => data <= "000000";
				when "000000100010011110" => data <= "000000";
				when "000000100010011111" => data <= "000000";
				when "000000101000000000" => data <= "000000";
				when "000000101000000001" => data <= "000000";
				when "000000101000000010" => data <= "000000";
				when "000000101000000011" => data <= "000000";
				when "000000101000000100" => data <= "000000";
				when "000000101000000101" => data <= "000000";
				when "000000101000000110" => data <= "000000";
				when "000000101000000111" => data <= "000000";
				when "000000101000001000" => data <= "000000";
				when "000000101000001001" => data <= "000000";
				when "000000101000001010" => data <= "000000";
				when "000000101000001011" => data <= "000000";
				when "000000101000001100" => data <= "000000";
				when "000000101000001101" => data <= "000000";
				when "000000101000001110" => data <= "000000";
				when "000000101000001111" => data <= "000000";
				when "000000101000010000" => data <= "000000";
				when "000000101000010001" => data <= "000000";
				when "000000101000010010" => data <= "000000";
				when "000000101000010011" => data <= "000000";
				when "000000101000010100" => data <= "000000";
				when "000000101000010101" => data <= "000000";
				when "000000101000010110" => data <= "000000";
				when "000000101000010111" => data <= "000000";
				when "000000101000011000" => data <= "000000";
				when "000000101000011001" => data <= "000000";
				when "000000101000011010" => data <= "000000";
				when "000000101000011011" => data <= "000000";
				when "000000101000011100" => data <= "000000";
				when "000000101000011101" => data <= "000000";
				when "000000101000011110" => data <= "000000";
				when "000000101000011111" => data <= "000000";
				when "000000101000100000" => data <= "000000";
				when "000000101000100001" => data <= "000000";
				when "000000101000100010" => data <= "000000";
				when "000000101000100011" => data <= "000000";
				when "000000101000100100" => data <= "000000";
				when "000000101000100101" => data <= "000000";
				when "000000101000100110" => data <= "000000";
				when "000000101000100111" => data <= "000000";
				when "000000101000101000" => data <= "000000";
				when "000000101000101001" => data <= "000000";
				when "000000101000101010" => data <= "000000";
				when "000000101000101011" => data <= "000000";
				when "000000101000101100" => data <= "000000";
				when "000000101000101101" => data <= "000000";
				when "000000101000101110" => data <= "000000";
				when "000000101000101111" => data <= "000000";
				when "000000101000110000" => data <= "000000";
				when "000000101000110001" => data <= "000000";
				when "000000101000110010" => data <= "000000";
				when "000000101000110011" => data <= "000000";
				when "000000101000110100" => data <= "000000";
				when "000000101000110101" => data <= "000000";
				when "000000101000110110" => data <= "000000";
				when "000000101000110111" => data <= "000000";
				when "000000101000111000" => data <= "000000";
				when "000000101000111001" => data <= "000000";
				when "000000101000111010" => data <= "000000";
				when "000000101000111011" => data <= "000000";
				when "000000101000111100" => data <= "000000";
				when "000000101000111101" => data <= "000000";
				when "000000101000111110" => data <= "000000";
				when "000000101000111111" => data <= "000000";
				when "000000101001000000" => data <= "000000";
				when "000000101001000001" => data <= "000000";
				when "000000101001000010" => data <= "000000";
				when "000000101001000011" => data <= "000000";
				when "000000101001000100" => data <= "000000";
				when "000000101001000101" => data <= "000000";
				when "000000101001000110" => data <= "000000";
				when "000000101001000111" => data <= "000000";
				when "000000101001001000" => data <= "000000";
				when "000000101001001001" => data <= "000000";
				when "000000101001001010" => data <= "000000";
				when "000000101001001011" => data <= "000000";
				when "000000101001001100" => data <= "000000";
				when "000000101001001101" => data <= "000000";
				when "000000101001001110" => data <= "000000";
				when "000000101001001111" => data <= "000000";
				when "000000101001010000" => data <= "000000";
				when "000000101001010001" => data <= "000000";
				when "000000101001010010" => data <= "000000";
				when "000000101001010011" => data <= "000000";
				when "000000101001010100" => data <= "000000";
				when "000000101001010101" => data <= "000000";
				when "000000101001010110" => data <= "000000";
				when "000000101001010111" => data <= "000000";
				when "000000101001011000" => data <= "000000";
				when "000000101001011001" => data <= "000000";
				when "000000101001011010" => data <= "000000";
				when "000000101001011011" => data <= "000000";
				when "000000101001011100" => data <= "000000";
				when "000000101001011101" => data <= "000000";
				when "000000101001011110" => data <= "000000";
				when "000000101001011111" => data <= "000000";
				when "000000101001100000" => data <= "000000";
				when "000000101001100001" => data <= "000000";
				when "000000101001100010" => data <= "000000";
				when "000000101001100011" => data <= "000000";
				when "000000101001100100" => data <= "000000";
				when "000000101001100101" => data <= "000000";
				when "000000101001100110" => data <= "000000";
				when "000000101001100111" => data <= "000000";
				when "000000101001101000" => data <= "000000";
				when "000000101001101001" => data <= "000000";
				when "000000101001101010" => data <= "000000";
				when "000000101001101011" => data <= "000000";
				when "000000101001101100" => data <= "000000";
				when "000000101001101101" => data <= "000000";
				when "000000101001101110" => data <= "000000";
				when "000000101001101111" => data <= "000000";
				when "000000101001110000" => data <= "000000";
				when "000000101001110001" => data <= "000000";
				when "000000101001110010" => data <= "000000";
				when "000000101001110011" => data <= "000000";
				when "000000101001110100" => data <= "000000";
				when "000000101001110101" => data <= "000000";
				when "000000101001110110" => data <= "000000";
				when "000000101001110111" => data <= "000000";
				when "000000101001111000" => data <= "000000";
				when "000000101001111001" => data <= "000000";
				when "000000101001111010" => data <= "000000";
				when "000000101001111011" => data <= "000000";
				when "000000101001111100" => data <= "000000";
				when "000000101001111101" => data <= "000000";
				when "000000101001111110" => data <= "000000";
				when "000000101001111111" => data <= "000000";
				when "000000101010000000" => data <= "000000";
				when "000000101010000001" => data <= "000000";
				when "000000101010000010" => data <= "000000";
				when "000000101010000011" => data <= "000000";
				when "000000101010000100" => data <= "000000";
				when "000000101010000101" => data <= "000000";
				when "000000101010000110" => data <= "000000";
				when "000000101010000111" => data <= "000000";
				when "000000101010001000" => data <= "000000";
				when "000000101010001001" => data <= "000000";
				when "000000101010001010" => data <= "000000";
				when "000000101010001011" => data <= "000000";
				when "000000101010001100" => data <= "000000";
				when "000000101010001101" => data <= "000000";
				when "000000101010001110" => data <= "000000";
				when "000000101010001111" => data <= "000000";
				when "000000101010010000" => data <= "000000";
				when "000000101010010001" => data <= "000000";
				when "000000101010010010" => data <= "000000";
				when "000000101010010011" => data <= "000000";
				when "000000101010010100" => data <= "000000";
				when "000000101010010101" => data <= "000000";
				when "000000101010010110" => data <= "000000";
				when "000000101010010111" => data <= "000000";
				when "000000101010011000" => data <= "000000";
				when "000000101010011001" => data <= "000000";
				when "000000101010011010" => data <= "000000";
				when "000000101010011011" => data <= "000000";
				when "000000101010011100" => data <= "000000";
				when "000000101010011101" => data <= "000000";
				when "000000101010011110" => data <= "000000";
				when "000000101010011111" => data <= "000000";
				when "000000110000000000" => data <= "000000";
				when "000000110000000001" => data <= "000000";
				when "000000110000000010" => data <= "000000";
				when "000000110000000011" => data <= "000000";
				when "000000110000000100" => data <= "000000";
				when "000000110000000101" => data <= "000000";
				when "000000110000000110" => data <= "000000";
				when "000000110000000111" => data <= "000000";
				when "000000110000001000" => data <= "000000";
				when "000000110000001001" => data <= "000000";
				when "000000110000001010" => data <= "000000";
				when "000000110000001011" => data <= "000000";
				when "000000110000001100" => data <= "000000";
				when "000000110000001101" => data <= "000000";
				when "000000110000001110" => data <= "000000";
				when "000000110000001111" => data <= "000000";
				when "000000110000010000" => data <= "000000";
				when "000000110000010001" => data <= "000000";
				when "000000110000010010" => data <= "000000";
				when "000000110000010011" => data <= "000000";
				when "000000110000010100" => data <= "000000";
				when "000000110000010101" => data <= "000000";
				when "000000110000010110" => data <= "000000";
				when "000000110000010111" => data <= "000000";
				when "000000110000011000" => data <= "000000";
				when "000000110000011001" => data <= "000000";
				when "000000110000011010" => data <= "000000";
				when "000000110000011011" => data <= "000000";
				when "000000110000011100" => data <= "000000";
				when "000000110000011101" => data <= "000000";
				when "000000110000011110" => data <= "000000";
				when "000000110000011111" => data <= "000000";
				when "000000110000100000" => data <= "000000";
				when "000000110000100001" => data <= "000000";
				when "000000110000100010" => data <= "000000";
				when "000000110000100011" => data <= "000000";
				when "000000110000100100" => data <= "000000";
				when "000000110000100101" => data <= "000000";
				when "000000110000100110" => data <= "000000";
				when "000000110000100111" => data <= "000000";
				when "000000110000101000" => data <= "000000";
				when "000000110000101001" => data <= "000000";
				when "000000110000101010" => data <= "000000";
				when "000000110000101011" => data <= "000000";
				when "000000110000101100" => data <= "000000";
				when "000000110000101101" => data <= "000000";
				when "000000110000101110" => data <= "000000";
				when "000000110000101111" => data <= "000000";
				when "000000110000110000" => data <= "000000";
				when "000000110000110001" => data <= "000000";
				when "000000110000110010" => data <= "000000";
				when "000000110000110011" => data <= "000000";
				when "000000110000110100" => data <= "000000";
				when "000000110000110101" => data <= "000000";
				when "000000110000110110" => data <= "000000";
				when "000000110000110111" => data <= "000000";
				when "000000110000111000" => data <= "000000";
				when "000000110000111001" => data <= "000000";
				when "000000110000111010" => data <= "000000";
				when "000000110000111011" => data <= "000000";
				when "000000110000111100" => data <= "000000";
				when "000000110000111101" => data <= "000000";
				when "000000110000111110" => data <= "000000";
				when "000000110000111111" => data <= "000000";
				when "000000110001000000" => data <= "000000";
				when "000000110001000001" => data <= "000000";
				when "000000110001000010" => data <= "000000";
				when "000000110001000011" => data <= "000000";
				when "000000110001000100" => data <= "000000";
				when "000000110001000101" => data <= "000000";
				when "000000110001000110" => data <= "000000";
				when "000000110001000111" => data <= "000000";
				when "000000110001001000" => data <= "000000";
				when "000000110001001001" => data <= "000000";
				when "000000110001001010" => data <= "000000";
				when "000000110001001011" => data <= "000000";
				when "000000110001001100" => data <= "000000";
				when "000000110001001101" => data <= "000000";
				when "000000110001001110" => data <= "000000";
				when "000000110001001111" => data <= "000000";
				when "000000110001010000" => data <= "000000";
				when "000000110001010001" => data <= "000000";
				when "000000110001010010" => data <= "000000";
				when "000000110001010011" => data <= "000000";
				when "000000110001010100" => data <= "000000";
				when "000000110001010101" => data <= "000000";
				when "000000110001010110" => data <= "000000";
				when "000000110001010111" => data <= "000000";
				when "000000110001011000" => data <= "000000";
				when "000000110001011001" => data <= "000000";
				when "000000110001011010" => data <= "000000";
				when "000000110001011011" => data <= "000000";
				when "000000110001011100" => data <= "000000";
				when "000000110001011101" => data <= "000000";
				when "000000110001011110" => data <= "000000";
				when "000000110001011111" => data <= "000000";
				when "000000110001100000" => data <= "000000";
				when "000000110001100001" => data <= "000000";
				when "000000110001100010" => data <= "000000";
				when "000000110001100011" => data <= "000000";
				when "000000110001100100" => data <= "000000";
				when "000000110001100101" => data <= "000000";
				when "000000110001100110" => data <= "000000";
				when "000000110001100111" => data <= "000000";
				when "000000110001101000" => data <= "000000";
				when "000000110001101001" => data <= "000000";
				when "000000110001101010" => data <= "000000";
				when "000000110001101011" => data <= "000000";
				when "000000110001101100" => data <= "000000";
				when "000000110001101101" => data <= "000000";
				when "000000110001101110" => data <= "000000";
				when "000000110001101111" => data <= "000000";
				when "000000110001110000" => data <= "000000";
				when "000000110001110001" => data <= "000000";
				when "000000110001110010" => data <= "000000";
				when "000000110001110011" => data <= "000000";
				when "000000110001110100" => data <= "000000";
				when "000000110001110101" => data <= "000000";
				when "000000110001110110" => data <= "000000";
				when "000000110001110111" => data <= "000000";
				when "000000110001111000" => data <= "000000";
				when "000000110001111001" => data <= "000000";
				when "000000110001111010" => data <= "000000";
				when "000000110001111011" => data <= "000000";
				when "000000110001111100" => data <= "000000";
				when "000000110001111101" => data <= "000000";
				when "000000110001111110" => data <= "000000";
				when "000000110001111111" => data <= "000000";
				when "000000110010000000" => data <= "000000";
				when "000000110010000001" => data <= "000000";
				when "000000110010000010" => data <= "000000";
				when "000000110010000011" => data <= "000000";
				when "000000110010000100" => data <= "000000";
				when "000000110010000101" => data <= "000000";
				when "000000110010000110" => data <= "000000";
				when "000000110010000111" => data <= "000000";
				when "000000110010001000" => data <= "000000";
				when "000000110010001001" => data <= "000000";
				when "000000110010001010" => data <= "000000";
				when "000000110010001011" => data <= "000000";
				when "000000110010001100" => data <= "000000";
				when "000000110010001101" => data <= "000000";
				when "000000110010001110" => data <= "000000";
				when "000000110010001111" => data <= "000000";
				when "000000110010010000" => data <= "000000";
				when "000000110010010001" => data <= "000000";
				when "000000110010010010" => data <= "000000";
				when "000000110010010011" => data <= "000000";
				when "000000110010010100" => data <= "000000";
				when "000000110010010101" => data <= "000000";
				when "000000110010010110" => data <= "000000";
				when "000000110010010111" => data <= "000000";
				when "000000110010011000" => data <= "000000";
				when "000000110010011001" => data <= "000000";
				when "000000110010011010" => data <= "000000";
				when "000000110010011011" => data <= "000000";
				when "000000110010011100" => data <= "000000";
				when "000000110010011101" => data <= "000000";
				when "000000110010011110" => data <= "000000";
				when "000000110010011111" => data <= "000000";
				when "000000111000000000" => data <= "000000";
				when "000000111000000001" => data <= "000000";
				when "000000111000000010" => data <= "000000";
				when "000000111000000011" => data <= "000000";
				when "000000111000000100" => data <= "000000";
				when "000000111000000101" => data <= "000000";
				when "000000111000000110" => data <= "000000";
				when "000000111000000111" => data <= "000000";
				when "000000111000001000" => data <= "000000";
				when "000000111000001001" => data <= "000000";
				when "000000111000001010" => data <= "000000";
				when "000000111000001011" => data <= "000000";
				when "000000111000001100" => data <= "000000";
				when "000000111000001101" => data <= "000000";
				when "000000111000001110" => data <= "000000";
				when "000000111000001111" => data <= "000000";
				when "000000111000010000" => data <= "000000";
				when "000000111000010001" => data <= "000000";
				when "000000111000010010" => data <= "000000";
				when "000000111000010011" => data <= "000000";
				when "000000111000010100" => data <= "000000";
				when "000000111000010101" => data <= "000000";
				when "000000111000010110" => data <= "000000";
				when "000000111000010111" => data <= "000000";
				when "000000111000011000" => data <= "000000";
				when "000000111000011001" => data <= "000000";
				when "000000111000011010" => data <= "000000";
				when "000000111000011011" => data <= "000000";
				when "000000111000011100" => data <= "000000";
				when "000000111000011101" => data <= "000000";
				when "000000111000011110" => data <= "000000";
				when "000000111000011111" => data <= "000000";
				when "000000111000100000" => data <= "000000";
				when "000000111000100001" => data <= "000000";
				when "000000111000100010" => data <= "000000";
				when "000000111000100011" => data <= "000000";
				when "000000111000100100" => data <= "000000";
				when "000000111000100101" => data <= "000000";
				when "000000111000100110" => data <= "000000";
				when "000000111000100111" => data <= "000000";
				when "000000111000101000" => data <= "000000";
				when "000000111000101001" => data <= "000000";
				when "000000111000101010" => data <= "000000";
				when "000000111000101011" => data <= "000000";
				when "000000111000101100" => data <= "000000";
				when "000000111000101101" => data <= "000000";
				when "000000111000101110" => data <= "000000";
				when "000000111000101111" => data <= "000000";
				when "000000111000110000" => data <= "000000";
				when "000000111000110001" => data <= "000000";
				when "000000111000110010" => data <= "000000";
				when "000000111000110011" => data <= "000000";
				when "000000111000110100" => data <= "000000";
				when "000000111000110101" => data <= "000000";
				when "000000111000110110" => data <= "000000";
				when "000000111000110111" => data <= "000000";
				when "000000111000111000" => data <= "000000";
				when "000000111000111001" => data <= "000000";
				when "000000111000111010" => data <= "000000";
				when "000000111000111011" => data <= "000000";
				when "000000111000111100" => data <= "000000";
				when "000000111000111101" => data <= "000000";
				when "000000111000111110" => data <= "000000";
				when "000000111000111111" => data <= "000000";
				when "000000111001000000" => data <= "000000";
				when "000000111001000001" => data <= "000000";
				when "000000111001000010" => data <= "000000";
				when "000000111001000011" => data <= "000000";
				when "000000111001000100" => data <= "000000";
				when "000000111001000101" => data <= "000000";
				when "000000111001000110" => data <= "000000";
				when "000000111001000111" => data <= "000000";
				when "000000111001001000" => data <= "000000";
				when "000000111001001001" => data <= "000000";
				when "000000111001001010" => data <= "000000";
				when "000000111001001011" => data <= "000000";
				when "000000111001001100" => data <= "000000";
				when "000000111001001101" => data <= "000000";
				when "000000111001001110" => data <= "000000";
				when "000000111001001111" => data <= "000000";
				when "000000111001010000" => data <= "000000";
				when "000000111001010001" => data <= "000000";
				when "000000111001010010" => data <= "000000";
				when "000000111001010011" => data <= "000000";
				when "000000111001010100" => data <= "000000";
				when "000000111001010101" => data <= "000000";
				when "000000111001010110" => data <= "000000";
				when "000000111001010111" => data <= "000000";
				when "000000111001011000" => data <= "000000";
				when "000000111001011001" => data <= "000000";
				when "000000111001011010" => data <= "000000";
				when "000000111001011011" => data <= "000000";
				when "000000111001011100" => data <= "000000";
				when "000000111001011101" => data <= "000000";
				when "000000111001011110" => data <= "000000";
				when "000000111001011111" => data <= "000000";
				when "000000111001100000" => data <= "000000";
				when "000000111001100001" => data <= "000000";
				when "000000111001100010" => data <= "000000";
				when "000000111001100011" => data <= "000000";
				when "000000111001100100" => data <= "000000";
				when "000000111001100101" => data <= "000000";
				when "000000111001100110" => data <= "000000";
				when "000000111001100111" => data <= "000000";
				when "000000111001101000" => data <= "000000";
				when "000000111001101001" => data <= "000000";
				when "000000111001101010" => data <= "000000";
				when "000000111001101011" => data <= "000000";
				when "000000111001101100" => data <= "000000";
				when "000000111001101101" => data <= "000000";
				when "000000111001101110" => data <= "000000";
				when "000000111001101111" => data <= "000000";
				when "000000111001110000" => data <= "000000";
				when "000000111001110001" => data <= "000000";
				when "000000111001110010" => data <= "000000";
				when "000000111001110011" => data <= "000000";
				when "000000111001110100" => data <= "000000";
				when "000000111001110101" => data <= "000000";
				when "000000111001110110" => data <= "000000";
				when "000000111001110111" => data <= "000000";
				when "000000111001111000" => data <= "000000";
				when "000000111001111001" => data <= "000000";
				when "000000111001111010" => data <= "000000";
				when "000000111001111011" => data <= "000000";
				when "000000111001111100" => data <= "000000";
				when "000000111001111101" => data <= "000000";
				when "000000111001111110" => data <= "000000";
				when "000000111001111111" => data <= "000000";
				when "000000111010000000" => data <= "000000";
				when "000000111010000001" => data <= "000000";
				when "000000111010000010" => data <= "000000";
				when "000000111010000011" => data <= "000000";
				when "000000111010000100" => data <= "000000";
				when "000000111010000101" => data <= "000000";
				when "000000111010000110" => data <= "000000";
				when "000000111010000111" => data <= "000000";
				when "000000111010001000" => data <= "000000";
				when "000000111010001001" => data <= "000000";
				when "000000111010001010" => data <= "000000";
				when "000000111010001011" => data <= "000000";
				when "000000111010001100" => data <= "000000";
				when "000000111010001101" => data <= "000000";
				when "000000111010001110" => data <= "000000";
				when "000000111010001111" => data <= "000000";
				when "000000111010010000" => data <= "000000";
				when "000000111010010001" => data <= "000000";
				when "000000111010010010" => data <= "000000";
				when "000000111010010011" => data <= "000000";
				when "000000111010010100" => data <= "000000";
				when "000000111010010101" => data <= "000000";
				when "000000111010010110" => data <= "000000";
				when "000000111010010111" => data <= "000000";
				when "000000111010011000" => data <= "000000";
				when "000000111010011001" => data <= "000000";
				when "000000111010011010" => data <= "000000";
				when "000000111010011011" => data <= "000000";
				when "000000111010011100" => data <= "000000";
				when "000000111010011101" => data <= "000000";
				when "000000111010011110" => data <= "000000";
				when "000000111010011111" => data <= "000000";
				when "000001000000000000" => data <= "000000";
				when "000001000000000001" => data <= "000000";
				when "000001000000000010" => data <= "000000";
				when "000001000000000011" => data <= "000000";
				when "000001000000000100" => data <= "000000";
				when "000001000000000101" => data <= "000000";
				when "000001000000000110" => data <= "000000";
				when "000001000000000111" => data <= "000000";
				when "000001000000001000" => data <= "000000";
				when "000001000000001001" => data <= "000000";
				when "000001000000001010" => data <= "000000";
				when "000001000000001011" => data <= "000000";
				when "000001000000001100" => data <= "000000";
				when "000001000000001101" => data <= "000000";
				when "000001000000001110" => data <= "000000";
				when "000001000000001111" => data <= "000000";
				when "000001000000010000" => data <= "000000";
				when "000001000000010001" => data <= "000000";
				when "000001000000010010" => data <= "000000";
				when "000001000000010011" => data <= "000000";
				when "000001000000010100" => data <= "000000";
				when "000001000000010101" => data <= "000000";
				when "000001000000010110" => data <= "000000";
				when "000001000000010111" => data <= "000000";
				when "000001000000011000" => data <= "000000";
				when "000001000000011001" => data <= "000000";
				when "000001000000011010" => data <= "000000";
				when "000001000000011011" => data <= "000000";
				when "000001000000011100" => data <= "000000";
				when "000001000000011101" => data <= "000000";
				when "000001000000011110" => data <= "000000";
				when "000001000000011111" => data <= "000000";
				when "000001000000100000" => data <= "000000";
				when "000001000000100001" => data <= "000000";
				when "000001000000100010" => data <= "000000";
				when "000001000000100011" => data <= "000000";
				when "000001000000100100" => data <= "000000";
				when "000001000000100101" => data <= "000000";
				when "000001000000100110" => data <= "000000";
				when "000001000000100111" => data <= "000000";
				when "000001000000101000" => data <= "000000";
				when "000001000000101001" => data <= "000000";
				when "000001000000101010" => data <= "000000";
				when "000001000000101011" => data <= "000000";
				when "000001000000101100" => data <= "000000";
				when "000001000000101101" => data <= "000000";
				when "000001000000101110" => data <= "000000";
				when "000001000000101111" => data <= "000000";
				when "000001000000110000" => data <= "000000";
				when "000001000000110001" => data <= "000000";
				when "000001000000110010" => data <= "000000";
				when "000001000000110011" => data <= "000000";
				when "000001000000110100" => data <= "000000";
				when "000001000000110101" => data <= "000000";
				when "000001000000110110" => data <= "000000";
				when "000001000000110111" => data <= "000000";
				when "000001000000111000" => data <= "000000";
				when "000001000000111001" => data <= "000000";
				when "000001000000111010" => data <= "000000";
				when "000001000000111011" => data <= "000000";
				when "000001000000111100" => data <= "000000";
				when "000001000000111101" => data <= "000000";
				when "000001000000111110" => data <= "000000";
				when "000001000000111111" => data <= "000000";
				when "000001000001000000" => data <= "000000";
				when "000001000001000001" => data <= "000000";
				when "000001000001000010" => data <= "000000";
				when "000001000001000011" => data <= "000000";
				when "000001000001000100" => data <= "000000";
				when "000001000001000101" => data <= "000000";
				when "000001000001000110" => data <= "000000";
				when "000001000001000111" => data <= "000000";
				when "000001000001001000" => data <= "000000";
				when "000001000001001001" => data <= "000000";
				when "000001000001001010" => data <= "000000";
				when "000001000001001011" => data <= "000000";
				when "000001000001001100" => data <= "000000";
				when "000001000001001101" => data <= "000000";
				when "000001000001001110" => data <= "000000";
				when "000001000001001111" => data <= "000000";
				when "000001000001010000" => data <= "000000";
				when "000001000001010001" => data <= "000000";
				when "000001000001010010" => data <= "000000";
				when "000001000001010011" => data <= "000000";
				when "000001000001010100" => data <= "000000";
				when "000001000001010101" => data <= "000000";
				when "000001000001010110" => data <= "000000";
				when "000001000001010111" => data <= "000000";
				when "000001000001011000" => data <= "000000";
				when "000001000001011001" => data <= "000000";
				when "000001000001011010" => data <= "000000";
				when "000001000001011011" => data <= "000000";
				when "000001000001011100" => data <= "000000";
				when "000001000001011101" => data <= "000000";
				when "000001000001011110" => data <= "000000";
				when "000001000001011111" => data <= "000000";
				when "000001000001100000" => data <= "000000";
				when "000001000001100001" => data <= "000000";
				when "000001000001100010" => data <= "000000";
				when "000001000001100011" => data <= "000000";
				when "000001000001100100" => data <= "000000";
				when "000001000001100101" => data <= "000000";
				when "000001000001100110" => data <= "000000";
				when "000001000001100111" => data <= "000000";
				when "000001000001101000" => data <= "000000";
				when "000001000001101001" => data <= "000000";
				when "000001000001101010" => data <= "000000";
				when "000001000001101011" => data <= "000000";
				when "000001000001101100" => data <= "000000";
				when "000001000001101101" => data <= "000000";
				when "000001000001101110" => data <= "000000";
				when "000001000001101111" => data <= "000000";
				when "000001000001110000" => data <= "000000";
				when "000001000001110001" => data <= "000000";
				when "000001000001110010" => data <= "000000";
				when "000001000001110011" => data <= "000000";
				when "000001000001110100" => data <= "000000";
				when "000001000001110101" => data <= "000000";
				when "000001000001110110" => data <= "000000";
				when "000001000001110111" => data <= "000000";
				when "000001000001111000" => data <= "000000";
				when "000001000001111001" => data <= "000000";
				when "000001000001111010" => data <= "000000";
				when "000001000001111011" => data <= "000000";
				when "000001000001111100" => data <= "000000";
				when "000001000001111101" => data <= "000000";
				when "000001000001111110" => data <= "000000";
				when "000001000001111111" => data <= "000000";
				when "000001000010000000" => data <= "000000";
				when "000001000010000001" => data <= "000000";
				when "000001000010000010" => data <= "000000";
				when "000001000010000011" => data <= "000000";
				when "000001000010000100" => data <= "000000";
				when "000001000010000101" => data <= "000000";
				when "000001000010000110" => data <= "000000";
				when "000001000010000111" => data <= "000000";
				when "000001000010001000" => data <= "000000";
				when "000001000010001001" => data <= "000000";
				when "000001000010001010" => data <= "000000";
				when "000001000010001011" => data <= "000000";
				when "000001000010001100" => data <= "000000";
				when "000001000010001101" => data <= "000000";
				when "000001000010001110" => data <= "000000";
				when "000001000010001111" => data <= "000000";
				when "000001000010010000" => data <= "000000";
				when "000001000010010001" => data <= "000000";
				when "000001000010010010" => data <= "000000";
				when "000001000010010011" => data <= "000000";
				when "000001000010010100" => data <= "000000";
				when "000001000010010101" => data <= "000000";
				when "000001000010010110" => data <= "000000";
				when "000001000010010111" => data <= "000000";
				when "000001000010011000" => data <= "000000";
				when "000001000010011001" => data <= "000000";
				when "000001000010011010" => data <= "000000";
				when "000001000010011011" => data <= "000000";
				when "000001000010011100" => data <= "000000";
				when "000001000010011101" => data <= "000000";
				when "000001000010011110" => data <= "000000";
				when "000001000010011111" => data <= "000000";
				when "000001001000000000" => data <= "000000";
				when "000001001000000001" => data <= "000000";
				when "000001001000000010" => data <= "000000";
				when "000001001000000011" => data <= "000000";
				when "000001001000000100" => data <= "000000";
				when "000001001000000101" => data <= "000000";
				when "000001001000000110" => data <= "000000";
				when "000001001000000111" => data <= "000000";
				when "000001001000001000" => data <= "000000";
				when "000001001000001001" => data <= "000000";
				when "000001001000001010" => data <= "000000";
				when "000001001000001011" => data <= "000000";
				when "000001001000001100" => data <= "000000";
				when "000001001000001101" => data <= "000000";
				when "000001001000001110" => data <= "000000";
				when "000001001000001111" => data <= "000000";
				when "000001001000010000" => data <= "000000";
				when "000001001000010001" => data <= "000000";
				when "000001001000010010" => data <= "000000";
				when "000001001000010011" => data <= "000000";
				when "000001001000010100" => data <= "000000";
				when "000001001000010101" => data <= "000000";
				when "000001001000010110" => data <= "000000";
				when "000001001000010111" => data <= "000000";
				when "000001001000011000" => data <= "000000";
				when "000001001000011001" => data <= "000000";
				when "000001001000011010" => data <= "000000";
				when "000001001000011011" => data <= "000000";
				when "000001001000011100" => data <= "000000";
				when "000001001000011101" => data <= "000000";
				when "000001001000011110" => data <= "000000";
				when "000001001000011111" => data <= "000000";
				when "000001001000100000" => data <= "000000";
				when "000001001000100001" => data <= "000000";
				when "000001001000100010" => data <= "000000";
				when "000001001000100011" => data <= "000000";
				when "000001001000100100" => data <= "000000";
				when "000001001000100101" => data <= "000000";
				when "000001001000100110" => data <= "000000";
				when "000001001000100111" => data <= "000000";
				when "000001001000101000" => data <= "000000";
				when "000001001000101001" => data <= "000000";
				when "000001001000101010" => data <= "000000";
				when "000001001000101011" => data <= "000000";
				when "000001001000101100" => data <= "000000";
				when "000001001000101101" => data <= "000000";
				when "000001001000101110" => data <= "000000";
				when "000001001000101111" => data <= "000000";
				when "000001001000110000" => data <= "000000";
				when "000001001000110001" => data <= "000000";
				when "000001001000110010" => data <= "000000";
				when "000001001000110011" => data <= "000000";
				when "000001001000110100" => data <= "000000";
				when "000001001000110101" => data <= "000000";
				when "000001001000110110" => data <= "000000";
				when "000001001000110111" => data <= "000000";
				when "000001001000111000" => data <= "000000";
				when "000001001000111001" => data <= "000000";
				when "000001001000111010" => data <= "000000";
				when "000001001000111011" => data <= "000000";
				when "000001001000111100" => data <= "000000";
				when "000001001000111101" => data <= "000000";
				when "000001001000111110" => data <= "000000";
				when "000001001000111111" => data <= "000000";
				when "000001001001000000" => data <= "000000";
				when "000001001001000001" => data <= "000000";
				when "000001001001000010" => data <= "000000";
				when "000001001001000011" => data <= "000000";
				when "000001001001000100" => data <= "000000";
				when "000001001001000101" => data <= "000000";
				when "000001001001000110" => data <= "000000";
				when "000001001001000111" => data <= "000000";
				when "000001001001001000" => data <= "000000";
				when "000001001001001001" => data <= "000000";
				when "000001001001001010" => data <= "000000";
				when "000001001001001011" => data <= "000000";
				when "000001001001001100" => data <= "000000";
				when "000001001001001101" => data <= "000000";
				when "000001001001001110" => data <= "000000";
				when "000001001001001111" => data <= "000000";
				when "000001001001010000" => data <= "000000";
				when "000001001001010001" => data <= "000000";
				when "000001001001010010" => data <= "000000";
				when "000001001001010011" => data <= "000000";
				when "000001001001010100" => data <= "000000";
				when "000001001001010101" => data <= "000000";
				when "000001001001010110" => data <= "000000";
				when "000001001001010111" => data <= "000000";
				when "000001001001011000" => data <= "000000";
				when "000001001001011001" => data <= "000000";
				when "000001001001011010" => data <= "000000";
				when "000001001001011011" => data <= "000000";
				when "000001001001011100" => data <= "000000";
				when "000001001001011101" => data <= "000000";
				when "000001001001011110" => data <= "000000";
				when "000001001001011111" => data <= "000000";
				when "000001001001100000" => data <= "000000";
				when "000001001001100001" => data <= "000000";
				when "000001001001100010" => data <= "000000";
				when "000001001001100011" => data <= "000000";
				when "000001001001100100" => data <= "000000";
				when "000001001001100101" => data <= "000000";
				when "000001001001100110" => data <= "000000";
				when "000001001001100111" => data <= "000000";
				when "000001001001101000" => data <= "000000";
				when "000001001001101001" => data <= "000000";
				when "000001001001101010" => data <= "000000";
				when "000001001001101011" => data <= "000000";
				when "000001001001101100" => data <= "000000";
				when "000001001001101101" => data <= "000000";
				when "000001001001101110" => data <= "000000";
				when "000001001001101111" => data <= "000000";
				when "000001001001110000" => data <= "000000";
				when "000001001001110001" => data <= "000000";
				when "000001001001110010" => data <= "000000";
				when "000001001001110011" => data <= "000000";
				when "000001001001110100" => data <= "000000";
				when "000001001001110101" => data <= "000000";
				when "000001001001110110" => data <= "000000";
				when "000001001001110111" => data <= "000000";
				when "000001001001111000" => data <= "000000";
				when "000001001001111001" => data <= "000000";
				when "000001001001111010" => data <= "000000";
				when "000001001001111011" => data <= "000000";
				when "000001001001111100" => data <= "000000";
				when "000001001001111101" => data <= "000000";
				when "000001001001111110" => data <= "000000";
				when "000001001001111111" => data <= "000000";
				when "000001001010000000" => data <= "000000";
				when "000001001010000001" => data <= "000000";
				when "000001001010000010" => data <= "000000";
				when "000001001010000011" => data <= "000000";
				when "000001001010000100" => data <= "000000";
				when "000001001010000101" => data <= "000000";
				when "000001001010000110" => data <= "000000";
				when "000001001010000111" => data <= "000000";
				when "000001001010001000" => data <= "000000";
				when "000001001010001001" => data <= "000000";
				when "000001001010001010" => data <= "000000";
				when "000001001010001011" => data <= "000000";
				when "000001001010001100" => data <= "000000";
				when "000001001010001101" => data <= "000000";
				when "000001001010001110" => data <= "000000";
				when "000001001010001111" => data <= "000000";
				when "000001001010010000" => data <= "000000";
				when "000001001010010001" => data <= "000000";
				when "000001001010010010" => data <= "000000";
				when "000001001010010011" => data <= "000000";
				when "000001001010010100" => data <= "000000";
				when "000001001010010101" => data <= "000000";
				when "000001001010010110" => data <= "000000";
				when "000001001010010111" => data <= "000000";
				when "000001001010011000" => data <= "000000";
				when "000001001010011001" => data <= "000000";
				when "000001001010011010" => data <= "000000";
				when "000001001010011011" => data <= "000000";
				when "000001001010011100" => data <= "000000";
				when "000001001010011101" => data <= "000000";
				when "000001001010011110" => data <= "000000";
				when "000001001010011111" => data <= "000000";
				when "000001010000000000" => data <= "000000";
				when "000001010000000001" => data <= "000000";
				when "000001010000000010" => data <= "000000";
				when "000001010000000011" => data <= "000000";
				when "000001010000000100" => data <= "000000";
				when "000001010000000101" => data <= "000000";
				when "000001010000000110" => data <= "000000";
				when "000001010000000111" => data <= "000000";
				when "000001010000001000" => data <= "000000";
				when "000001010000001001" => data <= "000000";
				when "000001010000001010" => data <= "000000";
				when "000001010000001011" => data <= "000000";
				when "000001010000001100" => data <= "000000";
				when "000001010000001101" => data <= "000000";
				when "000001010000001110" => data <= "000000";
				when "000001010000001111" => data <= "000000";
				when "000001010000010000" => data <= "000000";
				when "000001010000010001" => data <= "000000";
				when "000001010000010010" => data <= "000000";
				when "000001010000010011" => data <= "000000";
				when "000001010000010100" => data <= "000000";
				when "000001010000010101" => data <= "000000";
				when "000001010000010110" => data <= "000000";
				when "000001010000010111" => data <= "000000";
				when "000001010000011000" => data <= "000000";
				when "000001010000011001" => data <= "000000";
				when "000001010000011010" => data <= "000000";
				when "000001010000011011" => data <= "000000";
				when "000001010000011100" => data <= "000000";
				when "000001010000011101" => data <= "000000";
				when "000001010000011110" => data <= "000000";
				when "000001010000011111" => data <= "000000";
				when "000001010000100000" => data <= "000000";
				when "000001010000100001" => data <= "000000";
				when "000001010000100010" => data <= "000000";
				when "000001010000100011" => data <= "000000";
				when "000001010000100100" => data <= "000000";
				when "000001010000100101" => data <= "000000";
				when "000001010000100110" => data <= "000000";
				when "000001010000100111" => data <= "000000";
				when "000001010000101000" => data <= "000000";
				when "000001010000101001" => data <= "000000";
				when "000001010000101010" => data <= "000000";
				when "000001010000101011" => data <= "000000";
				when "000001010000101100" => data <= "000000";
				when "000001010000101101" => data <= "000000";
				when "000001010000101110" => data <= "000000";
				when "000001010000101111" => data <= "000000";
				when "000001010000110000" => data <= "000000";
				when "000001010000110001" => data <= "000000";
				when "000001010000110010" => data <= "000000";
				when "000001010000110011" => data <= "000000";
				when "000001010000110100" => data <= "000000";
				when "000001010000110101" => data <= "000000";
				when "000001010000110110" => data <= "000000";
				when "000001010000110111" => data <= "000000";
				when "000001010000111000" => data <= "000000";
				when "000001010000111001" => data <= "000000";
				when "000001010000111010" => data <= "000000";
				when "000001010000111011" => data <= "000000";
				when "000001010000111100" => data <= "000000";
				when "000001010000111101" => data <= "000000";
				when "000001010000111110" => data <= "000000";
				when "000001010000111111" => data <= "000000";
				when "000001010001000000" => data <= "000000";
				when "000001010001000001" => data <= "000000";
				when "000001010001000010" => data <= "000000";
				when "000001010001000011" => data <= "000000";
				when "000001010001000100" => data <= "000000";
				when "000001010001000101" => data <= "000000";
				when "000001010001000110" => data <= "000000";
				when "000001010001000111" => data <= "000000";
				when "000001010001001000" => data <= "000000";
				when "000001010001001001" => data <= "000000";
				when "000001010001001010" => data <= "000000";
				when "000001010001001011" => data <= "000000";
				when "000001010001001100" => data <= "000000";
				when "000001010001001101" => data <= "000000";
				when "000001010001001110" => data <= "000000";
				when "000001010001001111" => data <= "000000";
				when "000001010001010000" => data <= "000000";
				when "000001010001010001" => data <= "000000";
				when "000001010001010010" => data <= "000000";
				when "000001010001010011" => data <= "000000";
				when "000001010001010100" => data <= "000000";
				when "000001010001010101" => data <= "000000";
				when "000001010001010110" => data <= "000000";
				when "000001010001010111" => data <= "000000";
				when "000001010001011000" => data <= "000000";
				when "000001010001011001" => data <= "000000";
				when "000001010001011010" => data <= "000000";
				when "000001010001011011" => data <= "000000";
				when "000001010001011100" => data <= "000000";
				when "000001010001011101" => data <= "000000";
				when "000001010001011110" => data <= "000000";
				when "000001010001011111" => data <= "000000";
				when "000001010001100000" => data <= "000000";
				when "000001010001100001" => data <= "000000";
				when "000001010001100010" => data <= "000000";
				when "000001010001100011" => data <= "000000";
				when "000001010001100100" => data <= "000000";
				when "000001010001100101" => data <= "000000";
				when "000001010001100110" => data <= "000000";
				when "000001010001100111" => data <= "000000";
				when "000001010001101000" => data <= "000000";
				when "000001010001101001" => data <= "000000";
				when "000001010001101010" => data <= "000000";
				when "000001010001101011" => data <= "000000";
				when "000001010001101100" => data <= "000000";
				when "000001010001101101" => data <= "000000";
				when "000001010001101110" => data <= "000000";
				when "000001010001101111" => data <= "000000";
				when "000001010001110000" => data <= "000000";
				when "000001010001110001" => data <= "000000";
				when "000001010001110010" => data <= "000000";
				when "000001010001110011" => data <= "000000";
				when "000001010001110100" => data <= "000000";
				when "000001010001110101" => data <= "000000";
				when "000001010001110110" => data <= "000000";
				when "000001010001110111" => data <= "000000";
				when "000001010001111000" => data <= "000000";
				when "000001010001111001" => data <= "000000";
				when "000001010001111010" => data <= "000000";
				when "000001010001111011" => data <= "000000";
				when "000001010001111100" => data <= "000000";
				when "000001010001111101" => data <= "000000";
				when "000001010001111110" => data <= "000000";
				when "000001010001111111" => data <= "000000";
				when "000001010010000000" => data <= "000000";
				when "000001010010000001" => data <= "000000";
				when "000001010010000010" => data <= "000000";
				when "000001010010000011" => data <= "000000";
				when "000001010010000100" => data <= "000000";
				when "000001010010000101" => data <= "000000";
				when "000001010010000110" => data <= "000000";
				when "000001010010000111" => data <= "000000";
				when "000001010010001000" => data <= "000000";
				when "000001010010001001" => data <= "000000";
				when "000001010010001010" => data <= "000000";
				when "000001010010001011" => data <= "000000";
				when "000001010010001100" => data <= "000000";
				when "000001010010001101" => data <= "000000";
				when "000001010010001110" => data <= "000000";
				when "000001010010001111" => data <= "000000";
				when "000001010010010000" => data <= "000000";
				when "000001010010010001" => data <= "000000";
				when "000001010010010010" => data <= "000000";
				when "000001010010010011" => data <= "000000";
				when "000001010010010100" => data <= "000000";
				when "000001010010010101" => data <= "000000";
				when "000001010010010110" => data <= "000000";
				when "000001010010010111" => data <= "000000";
				when "000001010010011000" => data <= "000000";
				when "000001010010011001" => data <= "000000";
				when "000001010010011010" => data <= "000000";
				when "000001010010011011" => data <= "000000";
				when "000001010010011100" => data <= "000000";
				when "000001010010011101" => data <= "000000";
				when "000001010010011110" => data <= "000000";
				when "000001010010011111" => data <= "000000";
				when "000001011000000000" => data <= "000000";
				when "000001011000000001" => data <= "000000";
				when "000001011000000010" => data <= "000000";
				when "000001011000000011" => data <= "000000";
				when "000001011000000100" => data <= "000000";
				when "000001011000000101" => data <= "000000";
				when "000001011000000110" => data <= "000000";
				when "000001011000000111" => data <= "000000";
				when "000001011000001000" => data <= "000000";
				when "000001011000001001" => data <= "000000";
				when "000001011000001010" => data <= "000000";
				when "000001011000001011" => data <= "000000";
				when "000001011000001100" => data <= "000000";
				when "000001011000001101" => data <= "000000";
				when "000001011000001110" => data <= "000000";
				when "000001011000001111" => data <= "000000";
				when "000001011000010000" => data <= "000000";
				when "000001011000010001" => data <= "000000";
				when "000001011000010010" => data <= "000000";
				when "000001011000010011" => data <= "000000";
				when "000001011000010100" => data <= "000000";
				when "000001011000010101" => data <= "000000";
				when "000001011000010110" => data <= "000000";
				when "000001011000010111" => data <= "000000";
				when "000001011000011000" => data <= "000000";
				when "000001011000011001" => data <= "000000";
				when "000001011000011010" => data <= "000000";
				when "000001011000011011" => data <= "000000";
				when "000001011000011100" => data <= "000000";
				when "000001011000011101" => data <= "000000";
				when "000001011000011110" => data <= "000000";
				when "000001011000011111" => data <= "000000";
				when "000001011000100000" => data <= "000000";
				when "000001011000100001" => data <= "000000";
				when "000001011000100010" => data <= "000000";
				when "000001011000100011" => data <= "000000";
				when "000001011000100100" => data <= "000000";
				when "000001011000100101" => data <= "000000";
				when "000001011000100110" => data <= "000000";
				when "000001011000100111" => data <= "000000";
				when "000001011000101000" => data <= "000000";
				when "000001011000101001" => data <= "000000";
				when "000001011000101010" => data <= "000000";
				when "000001011000101011" => data <= "000000";
				when "000001011000101100" => data <= "000000";
				when "000001011000101101" => data <= "000000";
				when "000001011000101110" => data <= "000000";
				when "000001011000101111" => data <= "000000";
				when "000001011000110000" => data <= "000000";
				when "000001011000110001" => data <= "000000";
				when "000001011000110010" => data <= "000000";
				when "000001011000110011" => data <= "000000";
				when "000001011000110100" => data <= "000000";
				when "000001011000110101" => data <= "000000";
				when "000001011000110110" => data <= "000000";
				when "000001011000110111" => data <= "000000";
				when "000001011000111000" => data <= "000000";
				when "000001011000111001" => data <= "000000";
				when "000001011000111010" => data <= "000000";
				when "000001011000111011" => data <= "000000";
				when "000001011000111100" => data <= "000000";
				when "000001011000111101" => data <= "000000";
				when "000001011000111110" => data <= "000000";
				when "000001011000111111" => data <= "000000";
				when "000001011001000000" => data <= "000000";
				when "000001011001000001" => data <= "000000";
				when "000001011001000010" => data <= "000000";
				when "000001011001000011" => data <= "000000";
				when "000001011001000100" => data <= "000000";
				when "000001011001000101" => data <= "000000";
				when "000001011001000110" => data <= "000000";
				when "000001011001000111" => data <= "000000";
				when "000001011001001000" => data <= "000000";
				when "000001011001001001" => data <= "000000";
				when "000001011001001010" => data <= "000000";
				when "000001011001001011" => data <= "000000";
				when "000001011001001100" => data <= "000000";
				when "000001011001001101" => data <= "000000";
				when "000001011001001110" => data <= "000000";
				when "000001011001001111" => data <= "000000";
				when "000001011001010000" => data <= "000000";
				when "000001011001010001" => data <= "000000";
				when "000001011001010010" => data <= "000000";
				when "000001011001010011" => data <= "000000";
				when "000001011001010100" => data <= "000000";
				when "000001011001010101" => data <= "000000";
				when "000001011001010110" => data <= "000000";
				when "000001011001010111" => data <= "000000";
				when "000001011001011000" => data <= "000000";
				when "000001011001011001" => data <= "000000";
				when "000001011001011010" => data <= "000000";
				when "000001011001011011" => data <= "000000";
				when "000001011001011100" => data <= "000000";
				when "000001011001011101" => data <= "000000";
				when "000001011001011110" => data <= "000000";
				when "000001011001011111" => data <= "000000";
				when "000001011001100000" => data <= "000000";
				when "000001011001100001" => data <= "000000";
				when "000001011001100010" => data <= "000000";
				when "000001011001100011" => data <= "000000";
				when "000001011001100100" => data <= "000000";
				when "000001011001100101" => data <= "000000";
				when "000001011001100110" => data <= "000000";
				when "000001011001100111" => data <= "000000";
				when "000001011001101000" => data <= "000000";
				when "000001011001101001" => data <= "000000";
				when "000001011001101010" => data <= "000000";
				when "000001011001101011" => data <= "000000";
				when "000001011001101100" => data <= "000000";
				when "000001011001101101" => data <= "000000";
				when "000001011001101110" => data <= "000000";
				when "000001011001101111" => data <= "000000";
				when "000001011001110000" => data <= "000000";
				when "000001011001110001" => data <= "000000";
				when "000001011001110010" => data <= "000000";
				when "000001011001110011" => data <= "000000";
				when "000001011001110100" => data <= "000000";
				when "000001011001110101" => data <= "000000";
				when "000001011001110110" => data <= "000000";
				when "000001011001110111" => data <= "000000";
				when "000001011001111000" => data <= "000000";
				when "000001011001111001" => data <= "000000";
				when "000001011001111010" => data <= "000000";
				when "000001011001111011" => data <= "000000";
				when "000001011001111100" => data <= "000000";
				when "000001011001111101" => data <= "000000";
				when "000001011001111110" => data <= "000000";
				when "000001011001111111" => data <= "000000";
				when "000001011010000000" => data <= "000000";
				when "000001011010000001" => data <= "000000";
				when "000001011010000010" => data <= "000000";
				when "000001011010000011" => data <= "000000";
				when "000001011010000100" => data <= "000000";
				when "000001011010000101" => data <= "000000";
				when "000001011010000110" => data <= "000000";
				when "000001011010000111" => data <= "000000";
				when "000001011010001000" => data <= "000000";
				when "000001011010001001" => data <= "000000";
				when "000001011010001010" => data <= "000000";
				when "000001011010001011" => data <= "000000";
				when "000001011010001100" => data <= "000000";
				when "000001011010001101" => data <= "000000";
				when "000001011010001110" => data <= "000000";
				when "000001011010001111" => data <= "000000";
				when "000001011010010000" => data <= "000000";
				when "000001011010010001" => data <= "000000";
				when "000001011010010010" => data <= "000000";
				when "000001011010010011" => data <= "000000";
				when "000001011010010100" => data <= "000000";
				when "000001011010010101" => data <= "000000";
				when "000001011010010110" => data <= "000000";
				when "000001011010010111" => data <= "000000";
				when "000001011010011000" => data <= "000000";
				when "000001011010011001" => data <= "000000";
				when "000001011010011010" => data <= "000000";
				when "000001011010011011" => data <= "000000";
				when "000001011010011100" => data <= "000000";
				when "000001011010011101" => data <= "000000";
				when "000001011010011110" => data <= "000000";
				when "000001011010011111" => data <= "000000";
				when "000001100000000000" => data <= "000000";
				when "000001100000000001" => data <= "000000";
				when "000001100000000010" => data <= "000000";
				when "000001100000000011" => data <= "000000";
				when "000001100000000100" => data <= "000000";
				when "000001100000000101" => data <= "000000";
				when "000001100000000110" => data <= "000000";
				when "000001100000000111" => data <= "000000";
				when "000001100000001000" => data <= "000000";
				when "000001100000001001" => data <= "000000";
				when "000001100000001010" => data <= "000000";
				when "000001100000001011" => data <= "000000";
				when "000001100000001100" => data <= "000000";
				when "000001100000001101" => data <= "000000";
				when "000001100000001110" => data <= "000000";
				when "000001100000001111" => data <= "000000";
				when "000001100000010000" => data <= "000000";
				when "000001100000010001" => data <= "000000";
				when "000001100000010010" => data <= "000000";
				when "000001100000010011" => data <= "000000";
				when "000001100000010100" => data <= "000000";
				when "000001100000010101" => data <= "000000";
				when "000001100000010110" => data <= "000000";
				when "000001100000010111" => data <= "000000";
				when "000001100000011000" => data <= "000000";
				when "000001100000011001" => data <= "000000";
				when "000001100000011010" => data <= "000000";
				when "000001100000011011" => data <= "000000";
				when "000001100000011100" => data <= "000000";
				when "000001100000011101" => data <= "000000";
				when "000001100000011110" => data <= "000000";
				when "000001100000011111" => data <= "000000";
				when "000001100000100000" => data <= "000000";
				when "000001100000100001" => data <= "000000";
				when "000001100000100010" => data <= "000000";
				when "000001100000100011" => data <= "000000";
				when "000001100000100100" => data <= "000000";
				when "000001100000100101" => data <= "000000";
				when "000001100000100110" => data <= "000000";
				when "000001100000100111" => data <= "000000";
				when "000001100000101000" => data <= "000000";
				when "000001100000101001" => data <= "000000";
				when "000001100000101010" => data <= "000000";
				when "000001100000101011" => data <= "000000";
				when "000001100000101100" => data <= "000000";
				when "000001100000101101" => data <= "000000";
				when "000001100000101110" => data <= "000000";
				when "000001100000101111" => data <= "000000";
				when "000001100000110000" => data <= "000000";
				when "000001100000110001" => data <= "000000";
				when "000001100000110010" => data <= "000000";
				when "000001100000110011" => data <= "000000";
				when "000001100000110100" => data <= "000000";
				when "000001100000110101" => data <= "000000";
				when "000001100000110110" => data <= "000000";
				when "000001100000110111" => data <= "000000";
				when "000001100000111000" => data <= "000000";
				when "000001100000111001" => data <= "000000";
				when "000001100000111010" => data <= "000000";
				when "000001100000111011" => data <= "000000";
				when "000001100000111100" => data <= "000000";
				when "000001100000111101" => data <= "000000";
				when "000001100000111110" => data <= "000000";
				when "000001100000111111" => data <= "000000";
				when "000001100001000000" => data <= "000000";
				when "000001100001000001" => data <= "000000";
				when "000001100001000010" => data <= "000000";
				when "000001100001000011" => data <= "000000";
				when "000001100001000100" => data <= "000000";
				when "000001100001000101" => data <= "000000";
				when "000001100001000110" => data <= "000000";
				when "000001100001000111" => data <= "000000";
				when "000001100001001000" => data <= "000000";
				when "000001100001001001" => data <= "000000";
				when "000001100001001010" => data <= "000000";
				when "000001100001001011" => data <= "000000";
				when "000001100001001100" => data <= "000000";
				when "000001100001001101" => data <= "000000";
				when "000001100001001110" => data <= "000000";
				when "000001100001001111" => data <= "000000";
				when "000001100001010000" => data <= "000000";
				when "000001100001010001" => data <= "000000";
				when "000001100001010010" => data <= "000000";
				when "000001100001010011" => data <= "000000";
				when "000001100001010100" => data <= "000000";
				when "000001100001010101" => data <= "000000";
				when "000001100001010110" => data <= "000000";
				when "000001100001010111" => data <= "000000";
				when "000001100001011000" => data <= "000000";
				when "000001100001011001" => data <= "000000";
				when "000001100001011010" => data <= "000000";
				when "000001100001011011" => data <= "000000";
				when "000001100001011100" => data <= "000000";
				when "000001100001011101" => data <= "000000";
				when "000001100001011110" => data <= "000000";
				when "000001100001011111" => data <= "000000";
				when "000001100001100000" => data <= "000000";
				when "000001100001100001" => data <= "000000";
				when "000001100001100010" => data <= "000000";
				when "000001100001100011" => data <= "000000";
				when "000001100001100100" => data <= "000000";
				when "000001100001100101" => data <= "000000";
				when "000001100001100110" => data <= "000000";
				when "000001100001100111" => data <= "000000";
				when "000001100001101000" => data <= "000000";
				when "000001100001101001" => data <= "000000";
				when "000001100001101010" => data <= "000000";
				when "000001100001101011" => data <= "000000";
				when "000001100001101100" => data <= "000000";
				when "000001100001101101" => data <= "000000";
				when "000001100001101110" => data <= "000000";
				when "000001100001101111" => data <= "000000";
				when "000001100001110000" => data <= "000000";
				when "000001100001110001" => data <= "000000";
				when "000001100001110010" => data <= "000000";
				when "000001100001110011" => data <= "000000";
				when "000001100001110100" => data <= "000000";
				when "000001100001110101" => data <= "000000";
				when "000001100001110110" => data <= "000000";
				when "000001100001110111" => data <= "000000";
				when "000001100001111000" => data <= "000000";
				when "000001100001111001" => data <= "000000";
				when "000001100001111010" => data <= "000000";
				when "000001100001111011" => data <= "000000";
				when "000001100001111100" => data <= "000000";
				when "000001100001111101" => data <= "000000";
				when "000001100001111110" => data <= "000000";
				when "000001100001111111" => data <= "000000";
				when "000001100010000000" => data <= "000000";
				when "000001100010000001" => data <= "000000";
				when "000001100010000010" => data <= "000000";
				when "000001100010000011" => data <= "000000";
				when "000001100010000100" => data <= "000000";
				when "000001100010000101" => data <= "000000";
				when "000001100010000110" => data <= "000000";
				when "000001100010000111" => data <= "000000";
				when "000001100010001000" => data <= "000000";
				when "000001100010001001" => data <= "000000";
				when "000001100010001010" => data <= "000000";
				when "000001100010001011" => data <= "000000";
				when "000001100010001100" => data <= "000000";
				when "000001100010001101" => data <= "000000";
				when "000001100010001110" => data <= "000000";
				when "000001100010001111" => data <= "000000";
				when "000001100010010000" => data <= "000000";
				when "000001100010010001" => data <= "000000";
				when "000001100010010010" => data <= "000000";
				when "000001100010010011" => data <= "000000";
				when "000001100010010100" => data <= "000000";
				when "000001100010010101" => data <= "000000";
				when "000001100010010110" => data <= "000000";
				when "000001100010010111" => data <= "000000";
				when "000001100010011000" => data <= "000000";
				when "000001100010011001" => data <= "000000";
				when "000001100010011010" => data <= "000000";
				when "000001100010011011" => data <= "000000";
				when "000001100010011100" => data <= "000000";
				when "000001100010011101" => data <= "000000";
				when "000001100010011110" => data <= "000000";
				when "000001100010011111" => data <= "000000";
				when "000001101000000000" => data <= "000000";
				when "000001101000000001" => data <= "000000";
				when "000001101000000010" => data <= "000000";
				when "000001101000000011" => data <= "000000";
				when "000001101000000100" => data <= "000000";
				when "000001101000000101" => data <= "000000";
				when "000001101000000110" => data <= "000000";
				when "000001101000000111" => data <= "000000";
				when "000001101000001000" => data <= "000000";
				when "000001101000001001" => data <= "000000";
				when "000001101000001010" => data <= "000000";
				when "000001101000001011" => data <= "000000";
				when "000001101000001100" => data <= "000000";
				when "000001101000001101" => data <= "000000";
				when "000001101000001110" => data <= "000000";
				when "000001101000001111" => data <= "000000";
				when "000001101000010000" => data <= "000000";
				when "000001101000010001" => data <= "000000";
				when "000001101000010010" => data <= "000000";
				when "000001101000010011" => data <= "000000";
				when "000001101000010100" => data <= "000000";
				when "000001101000010101" => data <= "000000";
				when "000001101000010110" => data <= "000000";
				when "000001101000010111" => data <= "000000";
				when "000001101000011000" => data <= "000000";
				when "000001101000011001" => data <= "000000";
				when "000001101000011010" => data <= "000000";
				when "000001101000011011" => data <= "000000";
				when "000001101000011100" => data <= "000000";
				when "000001101000011101" => data <= "000000";
				when "000001101000011110" => data <= "000000";
				when "000001101000011111" => data <= "000000";
				when "000001101000100000" => data <= "000000";
				when "000001101000100001" => data <= "000000";
				when "000001101000100010" => data <= "000000";
				when "000001101000100011" => data <= "000000";
				when "000001101000100100" => data <= "000000";
				when "000001101000100101" => data <= "000000";
				when "000001101000100110" => data <= "000000";
				when "000001101000100111" => data <= "000000";
				when "000001101000101000" => data <= "000000";
				when "000001101000101001" => data <= "000000";
				when "000001101000101010" => data <= "000000";
				when "000001101000101011" => data <= "000000";
				when "000001101000101100" => data <= "000000";
				when "000001101000101101" => data <= "000000";
				when "000001101000101110" => data <= "000000";
				when "000001101000101111" => data <= "000000";
				when "000001101000110000" => data <= "000000";
				when "000001101000110001" => data <= "000000";
				when "000001101000110010" => data <= "000000";
				when "000001101000110011" => data <= "000000";
				when "000001101000110100" => data <= "000000";
				when "000001101000110101" => data <= "000000";
				when "000001101000110110" => data <= "000000";
				when "000001101000110111" => data <= "000000";
				when "000001101000111000" => data <= "000000";
				when "000001101000111001" => data <= "000000";
				when "000001101000111010" => data <= "000000";
				when "000001101000111011" => data <= "000000";
				when "000001101000111100" => data <= "000000";
				when "000001101000111101" => data <= "000000";
				when "000001101000111110" => data <= "000000";
				when "000001101000111111" => data <= "000000";
				when "000001101001000000" => data <= "000000";
				when "000001101001000001" => data <= "000000";
				when "000001101001000010" => data <= "000000";
				when "000001101001000011" => data <= "000000";
				when "000001101001000100" => data <= "000000";
				when "000001101001000101" => data <= "000000";
				when "000001101001000110" => data <= "000000";
				when "000001101001000111" => data <= "000000";
				when "000001101001001000" => data <= "000000";
				when "000001101001001001" => data <= "000000";
				when "000001101001001010" => data <= "000000";
				when "000001101001001011" => data <= "000000";
				when "000001101001001100" => data <= "000000";
				when "000001101001001101" => data <= "000000";
				when "000001101001001110" => data <= "000000";
				when "000001101001001111" => data <= "000000";
				when "000001101001010000" => data <= "000000";
				when "000001101001010001" => data <= "000000";
				when "000001101001010010" => data <= "000000";
				when "000001101001010011" => data <= "000000";
				when "000001101001010100" => data <= "000000";
				when "000001101001010101" => data <= "000000";
				when "000001101001010110" => data <= "000000";
				when "000001101001010111" => data <= "000000";
				when "000001101001011000" => data <= "000000";
				when "000001101001011001" => data <= "000000";
				when "000001101001011010" => data <= "000000";
				when "000001101001011011" => data <= "000000";
				when "000001101001011100" => data <= "000000";
				when "000001101001011101" => data <= "000000";
				when "000001101001011110" => data <= "000000";
				when "000001101001011111" => data <= "000000";
				when "000001101001100000" => data <= "000000";
				when "000001101001100001" => data <= "000000";
				when "000001101001100010" => data <= "000000";
				when "000001101001100011" => data <= "000000";
				when "000001101001100100" => data <= "000000";
				when "000001101001100101" => data <= "000000";
				when "000001101001100110" => data <= "000000";
				when "000001101001100111" => data <= "000000";
				when "000001101001101000" => data <= "000000";
				when "000001101001101001" => data <= "000000";
				when "000001101001101010" => data <= "000000";
				when "000001101001101011" => data <= "000000";
				when "000001101001101100" => data <= "000000";
				when "000001101001101101" => data <= "000000";
				when "000001101001101110" => data <= "000000";
				when "000001101001101111" => data <= "000000";
				when "000001101001110000" => data <= "000000";
				when "000001101001110001" => data <= "000000";
				when "000001101001110010" => data <= "000000";
				when "000001101001110011" => data <= "000000";
				when "000001101001110100" => data <= "000000";
				when "000001101001110101" => data <= "000000";
				when "000001101001110110" => data <= "000000";
				when "000001101001110111" => data <= "000000";
				when "000001101001111000" => data <= "000000";
				when "000001101001111001" => data <= "000000";
				when "000001101001111010" => data <= "000000";
				when "000001101001111011" => data <= "000000";
				when "000001101001111100" => data <= "000000";
				when "000001101001111101" => data <= "000000";
				when "000001101001111110" => data <= "000000";
				when "000001101001111111" => data <= "000000";
				when "000001101010000000" => data <= "000000";
				when "000001101010000001" => data <= "000000";
				when "000001101010000010" => data <= "000000";
				when "000001101010000011" => data <= "000000";
				when "000001101010000100" => data <= "000000";
				when "000001101010000101" => data <= "000000";
				when "000001101010000110" => data <= "000000";
				when "000001101010000111" => data <= "000000";
				when "000001101010001000" => data <= "000000";
				when "000001101010001001" => data <= "000000";
				when "000001101010001010" => data <= "000000";
				when "000001101010001011" => data <= "000000";
				when "000001101010001100" => data <= "000000";
				when "000001101010001101" => data <= "000000";
				when "000001101010001110" => data <= "000000";
				when "000001101010001111" => data <= "000000";
				when "000001101010010000" => data <= "000000";
				when "000001101010010001" => data <= "000000";
				when "000001101010010010" => data <= "000000";
				when "000001101010010011" => data <= "000000";
				when "000001101010010100" => data <= "000000";
				when "000001101010010101" => data <= "000000";
				when "000001101010010110" => data <= "000000";
				when "000001101010010111" => data <= "000000";
				when "000001101010011000" => data <= "000000";
				when "000001101010011001" => data <= "000000";
				when "000001101010011010" => data <= "000000";
				when "000001101010011011" => data <= "000000";
				when "000001101010011100" => data <= "000000";
				when "000001101010011101" => data <= "000000";
				when "000001101010011110" => data <= "000000";
				when "000001101010011111" => data <= "000000";
				when "000001110000000000" => data <= "000000";
				when "000001110000000001" => data <= "000000";
				when "000001110000000010" => data <= "000000";
				when "000001110000000011" => data <= "000000";
				when "000001110000000100" => data <= "000000";
				when "000001110000000101" => data <= "000000";
				when "000001110000000110" => data <= "000000";
				when "000001110000000111" => data <= "000000";
				when "000001110000001000" => data <= "000000";
				when "000001110000001001" => data <= "000000";
				when "000001110000001010" => data <= "000000";
				when "000001110000001011" => data <= "000000";
				when "000001110000001100" => data <= "000000";
				when "000001110000001101" => data <= "000000";
				when "000001110000001110" => data <= "000000";
				when "000001110000001111" => data <= "000000";
				when "000001110000010000" => data <= "000000";
				when "000001110000010001" => data <= "000000";
				when "000001110000010010" => data <= "000000";
				when "000001110000010011" => data <= "000000";
				when "000001110000010100" => data <= "000000";
				when "000001110000010101" => data <= "000000";
				when "000001110000010110" => data <= "000000";
				when "000001110000010111" => data <= "000000";
				when "000001110000011000" => data <= "000000";
				when "000001110000011001" => data <= "000000";
				when "000001110000011010" => data <= "000000";
				when "000001110000011011" => data <= "000000";
				when "000001110000011100" => data <= "000000";
				when "000001110000011101" => data <= "000000";
				when "000001110000011110" => data <= "000000";
				when "000001110000011111" => data <= "000000";
				when "000001110000100000" => data <= "000000";
				when "000001110000100001" => data <= "000000";
				when "000001110000100010" => data <= "000000";
				when "000001110000100011" => data <= "000000";
				when "000001110000100100" => data <= "000000";
				when "000001110000100101" => data <= "000000";
				when "000001110000100110" => data <= "000000";
				when "000001110000100111" => data <= "000000";
				when "000001110000101000" => data <= "000000";
				when "000001110000101001" => data <= "000000";
				when "000001110000101010" => data <= "000000";
				when "000001110000101011" => data <= "000000";
				when "000001110000101100" => data <= "000000";
				when "000001110000101101" => data <= "000000";
				when "000001110000101110" => data <= "000000";
				when "000001110000101111" => data <= "000000";
				when "000001110000110000" => data <= "000000";
				when "000001110000110001" => data <= "000000";
				when "000001110000110010" => data <= "000000";
				when "000001110000110011" => data <= "000000";
				when "000001110000110100" => data <= "000000";
				when "000001110000110101" => data <= "000000";
				when "000001110000110110" => data <= "000000";
				when "000001110000110111" => data <= "000000";
				when "000001110000111000" => data <= "000000";
				when "000001110000111001" => data <= "000000";
				when "000001110000111010" => data <= "000000";
				when "000001110000111011" => data <= "000000";
				when "000001110000111100" => data <= "000000";
				when "000001110000111101" => data <= "000000";
				when "000001110000111110" => data <= "000000";
				when "000001110000111111" => data <= "000000";
				when "000001110001000000" => data <= "000000";
				when "000001110001000001" => data <= "000000";
				when "000001110001000010" => data <= "000000";
				when "000001110001000011" => data <= "000000";
				when "000001110001000100" => data <= "000000";
				when "000001110001000101" => data <= "000000";
				when "000001110001000110" => data <= "000000";
				when "000001110001000111" => data <= "000000";
				when "000001110001001000" => data <= "000000";
				when "000001110001001001" => data <= "000000";
				when "000001110001001010" => data <= "000000";
				when "000001110001001011" => data <= "000000";
				when "000001110001001100" => data <= "000000";
				when "000001110001001101" => data <= "000000";
				when "000001110001001110" => data <= "000000";
				when "000001110001001111" => data <= "000000";
				when "000001110001010000" => data <= "000000";
				when "000001110001010001" => data <= "000000";
				when "000001110001010010" => data <= "000000";
				when "000001110001010011" => data <= "000000";
				when "000001110001010100" => data <= "000000";
				when "000001110001010101" => data <= "000000";
				when "000001110001010110" => data <= "000000";
				when "000001110001010111" => data <= "000000";
				when "000001110001011000" => data <= "000000";
				when "000001110001011001" => data <= "000000";
				when "000001110001011010" => data <= "000000";
				when "000001110001011011" => data <= "000000";
				when "000001110001011100" => data <= "000000";
				when "000001110001011101" => data <= "000000";
				when "000001110001011110" => data <= "000000";
				when "000001110001011111" => data <= "000000";
				when "000001110001100000" => data <= "000000";
				when "000001110001100001" => data <= "000000";
				when "000001110001100010" => data <= "000000";
				when "000001110001100011" => data <= "000000";
				when "000001110001100100" => data <= "000000";
				when "000001110001100101" => data <= "000000";
				when "000001110001100110" => data <= "000000";
				when "000001110001100111" => data <= "000000";
				when "000001110001101000" => data <= "000000";
				when "000001110001101001" => data <= "000000";
				when "000001110001101010" => data <= "000000";
				when "000001110001101011" => data <= "000000";
				when "000001110001101100" => data <= "000000";
				when "000001110001101101" => data <= "000000";
				when "000001110001101110" => data <= "000000";
				when "000001110001101111" => data <= "000000";
				when "000001110001110000" => data <= "000000";
				when "000001110001110001" => data <= "000000";
				when "000001110001110010" => data <= "000000";
				when "000001110001110011" => data <= "000000";
				when "000001110001110100" => data <= "000000";
				when "000001110001110101" => data <= "000000";
				when "000001110001110110" => data <= "000000";
				when "000001110001110111" => data <= "000000";
				when "000001110001111000" => data <= "000000";
				when "000001110001111001" => data <= "000000";
				when "000001110001111010" => data <= "000000";
				when "000001110001111011" => data <= "000000";
				when "000001110001111100" => data <= "000000";
				when "000001110001111101" => data <= "000000";
				when "000001110001111110" => data <= "000000";
				when "000001110001111111" => data <= "000000";
				when "000001110010000000" => data <= "000000";
				when "000001110010000001" => data <= "000000";
				when "000001110010000010" => data <= "000000";
				when "000001110010000011" => data <= "000000";
				when "000001110010000100" => data <= "000000";
				when "000001110010000101" => data <= "000000";
				when "000001110010000110" => data <= "000000";
				when "000001110010000111" => data <= "000000";
				when "000001110010001000" => data <= "000000";
				when "000001110010001001" => data <= "000000";
				when "000001110010001010" => data <= "000000";
				when "000001110010001011" => data <= "000000";
				when "000001110010001100" => data <= "000000";
				when "000001110010001101" => data <= "000000";
				when "000001110010001110" => data <= "000000";
				when "000001110010001111" => data <= "000000";
				when "000001110010010000" => data <= "000000";
				when "000001110010010001" => data <= "000000";
				when "000001110010010010" => data <= "000000";
				when "000001110010010011" => data <= "000000";
				when "000001110010010100" => data <= "000000";
				when "000001110010010101" => data <= "000000";
				when "000001110010010110" => data <= "000000";
				when "000001110010010111" => data <= "000000";
				when "000001110010011000" => data <= "000000";
				when "000001110010011001" => data <= "000000";
				when "000001110010011010" => data <= "000000";
				when "000001110010011011" => data <= "000000";
				when "000001110010011100" => data <= "000000";
				when "000001110010011101" => data <= "000000";
				when "000001110010011110" => data <= "000000";
				when "000001110010011111" => data <= "000000";
				when "000001111000000000" => data <= "000000";
				when "000001111000000001" => data <= "000000";
				when "000001111000000010" => data <= "000000";
				when "000001111000000011" => data <= "000000";
				when "000001111000000100" => data <= "000000";
				when "000001111000000101" => data <= "000000";
				when "000001111000000110" => data <= "000000";
				when "000001111000000111" => data <= "000000";
				when "000001111000001000" => data <= "000000";
				when "000001111000001001" => data <= "000000";
				when "000001111000001010" => data <= "000000";
				when "000001111000001011" => data <= "000000";
				when "000001111000001100" => data <= "000000";
				when "000001111000001101" => data <= "000000";
				when "000001111000001110" => data <= "000000";
				when "000001111000001111" => data <= "000000";
				when "000001111000010000" => data <= "000000";
				when "000001111000010001" => data <= "000000";
				when "000001111000010010" => data <= "000000";
				when "000001111000010011" => data <= "000000";
				when "000001111000010100" => data <= "000000";
				when "000001111000010101" => data <= "000000";
				when "000001111000010110" => data <= "000000";
				when "000001111000010111" => data <= "000000";
				when "000001111000011000" => data <= "000000";
				when "000001111000011001" => data <= "000000";
				when "000001111000011010" => data <= "000000";
				when "000001111000011011" => data <= "000000";
				when "000001111000011100" => data <= "000000";
				when "000001111000011101" => data <= "000000";
				when "000001111000011110" => data <= "000000";
				when "000001111000011111" => data <= "000000";
				when "000001111000100000" => data <= "000000";
				when "000001111000100001" => data <= "000000";
				when "000001111000100010" => data <= "000000";
				when "000001111000100011" => data <= "000000";
				when "000001111000100100" => data <= "000000";
				when "000001111000100101" => data <= "000000";
				when "000001111000100110" => data <= "000000";
				when "000001111000100111" => data <= "000000";
				when "000001111000101000" => data <= "000000";
				when "000001111000101001" => data <= "000000";
				when "000001111000101010" => data <= "000000";
				when "000001111000101011" => data <= "000000";
				when "000001111000101100" => data <= "000000";
				when "000001111000101101" => data <= "000000";
				when "000001111000101110" => data <= "000000";
				when "000001111000101111" => data <= "000000";
				when "000001111000110000" => data <= "000000";
				when "000001111000110001" => data <= "000000";
				when "000001111000110010" => data <= "000000";
				when "000001111000110011" => data <= "000000";
				when "000001111000110100" => data <= "000000";
				when "000001111000110101" => data <= "000000";
				when "000001111000110110" => data <= "000000";
				when "000001111000110111" => data <= "000000";
				when "000001111000111000" => data <= "000000";
				when "000001111000111001" => data <= "000000";
				when "000001111000111010" => data <= "000000";
				when "000001111000111011" => data <= "000000";
				when "000001111000111100" => data <= "000000";
				when "000001111000111101" => data <= "000000";
				when "000001111000111110" => data <= "000000";
				when "000001111000111111" => data <= "000000";
				when "000001111001000000" => data <= "000000";
				when "000001111001000001" => data <= "000000";
				when "000001111001000010" => data <= "000000";
				when "000001111001000011" => data <= "000000";
				when "000001111001000100" => data <= "000000";
				when "000001111001000101" => data <= "000000";
				when "000001111001000110" => data <= "000000";
				when "000001111001000111" => data <= "000000";
				when "000001111001001000" => data <= "000000";
				when "000001111001001001" => data <= "000000";
				when "000001111001001010" => data <= "000000";
				when "000001111001001011" => data <= "000000";
				when "000001111001001100" => data <= "000000";
				when "000001111001001101" => data <= "000000";
				when "000001111001001110" => data <= "000000";
				when "000001111001001111" => data <= "000000";
				when "000001111001010000" => data <= "000000";
				when "000001111001010001" => data <= "000000";
				when "000001111001010010" => data <= "000000";
				when "000001111001010011" => data <= "000000";
				when "000001111001010100" => data <= "000000";
				when "000001111001010101" => data <= "000000";
				when "000001111001010110" => data <= "000000";
				when "000001111001010111" => data <= "000000";
				when "000001111001011000" => data <= "000000";
				when "000001111001011001" => data <= "000000";
				when "000001111001011010" => data <= "000000";
				when "000001111001011011" => data <= "000000";
				when "000001111001011100" => data <= "000000";
				when "000001111001011101" => data <= "000000";
				when "000001111001011110" => data <= "000000";
				when "000001111001011111" => data <= "000000";
				when "000001111001100000" => data <= "000000";
				when "000001111001100001" => data <= "000000";
				when "000001111001100010" => data <= "000000";
				when "000001111001100011" => data <= "000000";
				when "000001111001100100" => data <= "000000";
				when "000001111001100101" => data <= "000000";
				when "000001111001100110" => data <= "000000";
				when "000001111001100111" => data <= "000000";
				when "000001111001101000" => data <= "000000";
				when "000001111001101001" => data <= "000000";
				when "000001111001101010" => data <= "000000";
				when "000001111001101011" => data <= "000000";
				when "000001111001101100" => data <= "000000";
				when "000001111001101101" => data <= "000000";
				when "000001111001101110" => data <= "000000";
				when "000001111001101111" => data <= "000000";
				when "000001111001110000" => data <= "000000";
				when "000001111001110001" => data <= "000000";
				when "000001111001110010" => data <= "000000";
				when "000001111001110011" => data <= "000000";
				when "000001111001110100" => data <= "000000";
				when "000001111001110101" => data <= "000000";
				when "000001111001110110" => data <= "000000";
				when "000001111001110111" => data <= "000000";
				when "000001111001111000" => data <= "000000";
				when "000001111001111001" => data <= "000000";
				when "000001111001111010" => data <= "000000";
				when "000001111001111011" => data <= "000000";
				when "000001111001111100" => data <= "000000";
				when "000001111001111101" => data <= "000000";
				when "000001111001111110" => data <= "000000";
				when "000001111001111111" => data <= "000000";
				when "000001111010000000" => data <= "000000";
				when "000001111010000001" => data <= "000000";
				when "000001111010000010" => data <= "000000";
				when "000001111010000011" => data <= "000000";
				when "000001111010000100" => data <= "000000";
				when "000001111010000101" => data <= "000000";
				when "000001111010000110" => data <= "000000";
				when "000001111010000111" => data <= "000000";
				when "000001111010001000" => data <= "000000";
				when "000001111010001001" => data <= "000000";
				when "000001111010001010" => data <= "000000";
				when "000001111010001011" => data <= "000000";
				when "000001111010001100" => data <= "000000";
				when "000001111010001101" => data <= "000000";
				when "000001111010001110" => data <= "000000";
				when "000001111010001111" => data <= "000000";
				when "000001111010010000" => data <= "000000";
				when "000001111010010001" => data <= "000000";
				when "000001111010010010" => data <= "000000";
				when "000001111010010011" => data <= "000000";
				when "000001111010010100" => data <= "000000";
				when "000001111010010101" => data <= "000000";
				when "000001111010010110" => data <= "000000";
				when "000001111010010111" => data <= "000000";
				when "000001111010011000" => data <= "000000";
				when "000001111010011001" => data <= "000000";
				when "000001111010011010" => data <= "000000";
				when "000001111010011011" => data <= "000000";
				when "000001111010011100" => data <= "000000";
				when "000001111010011101" => data <= "000000";
				when "000001111010011110" => data <= "000000";
				when "000001111010011111" => data <= "000000";
				when "000010000000000000" => data <= "000000";
				when "000010000000000001" => data <= "000000";
				when "000010000000000010" => data <= "000000";
				when "000010000000000011" => data <= "000000";
				when "000010000000000100" => data <= "000000";
				when "000010000000000101" => data <= "000000";
				when "000010000000000110" => data <= "000000";
				when "000010000000000111" => data <= "000000";
				when "000010000000001000" => data <= "000000";
				when "000010000000001001" => data <= "000000";
				when "000010000000001010" => data <= "000000";
				when "000010000000001011" => data <= "000000";
				when "000010000000001100" => data <= "000000";
				when "000010000000001101" => data <= "000000";
				when "000010000000001110" => data <= "000000";
				when "000010000000001111" => data <= "000000";
				when "000010000000010000" => data <= "000000";
				when "000010000000010001" => data <= "000000";
				when "000010000000010010" => data <= "000000";
				when "000010000000010011" => data <= "000000";
				when "000010000000010100" => data <= "000000";
				when "000010000000010101" => data <= "000000";
				when "000010000000010110" => data <= "000000";
				when "000010000000010111" => data <= "000000";
				when "000010000000011000" => data <= "000000";
				when "000010000000011001" => data <= "000000";
				when "000010000000011010" => data <= "000000";
				when "000010000000011011" => data <= "000000";
				when "000010000000011100" => data <= "000000";
				when "000010000000011101" => data <= "000000";
				when "000010000000011110" => data <= "000000";
				when "000010000000011111" => data <= "000000";
				when "000010000000100000" => data <= "000000";
				when "000010000000100001" => data <= "000000";
				when "000010000000100010" => data <= "000000";
				when "000010000000100011" => data <= "000000";
				when "000010000000100100" => data <= "000000";
				when "000010000000100101" => data <= "000000";
				when "000010000000100110" => data <= "000000";
				when "000010000000100111" => data <= "000000";
				when "000010000000101000" => data <= "000000";
				when "000010000000101001" => data <= "000000";
				when "000010000000101010" => data <= "000000";
				when "000010000000101011" => data <= "000000";
				when "000010000000101100" => data <= "000000";
				when "000010000000101101" => data <= "000000";
				when "000010000000101110" => data <= "000000";
				when "000010000000101111" => data <= "000000";
				when "000010000000110000" => data <= "000000";
				when "000010000000110001" => data <= "000000";
				when "000010000000110010" => data <= "000000";
				when "000010000000110011" => data <= "000000";
				when "000010000000110100" => data <= "000000";
				when "000010000000110101" => data <= "000000";
				when "000010000000110110" => data <= "000000";
				when "000010000000110111" => data <= "000000";
				when "000010000000111000" => data <= "000000";
				when "000010000000111001" => data <= "000000";
				when "000010000000111010" => data <= "000000";
				when "000010000000111011" => data <= "000000";
				when "000010000000111100" => data <= "000000";
				when "000010000000111101" => data <= "000000";
				when "000010000000111110" => data <= "000000";
				when "000010000000111111" => data <= "000000";
				when "000010000001000000" => data <= "000000";
				when "000010000001000001" => data <= "000000";
				when "000010000001000010" => data <= "000000";
				when "000010000001000011" => data <= "000000";
				when "000010000001000100" => data <= "000000";
				when "000010000001000101" => data <= "000000";
				when "000010000001000110" => data <= "000000";
				when "000010000001000111" => data <= "000000";
				when "000010000001001000" => data <= "000000";
				when "000010000001001001" => data <= "000000";
				when "000010000001001010" => data <= "000000";
				when "000010000001001011" => data <= "000000";
				when "000010000001001100" => data <= "000000";
				when "000010000001001101" => data <= "000000";
				when "000010000001001110" => data <= "000000";
				when "000010000001001111" => data <= "000000";
				when "000010000001010000" => data <= "000000";
				when "000010000001010001" => data <= "000000";
				when "000010000001010010" => data <= "000000";
				when "000010000001010011" => data <= "000000";
				when "000010000001010100" => data <= "000000";
				when "000010000001010101" => data <= "000000";
				when "000010000001010110" => data <= "000000";
				when "000010000001010111" => data <= "000000";
				when "000010000001011000" => data <= "000000";
				when "000010000001011001" => data <= "000000";
				when "000010000001011010" => data <= "000000";
				when "000010000001011011" => data <= "000000";
				when "000010000001011100" => data <= "000000";
				when "000010000001011101" => data <= "000000";
				when "000010000001011110" => data <= "000000";
				when "000010000001011111" => data <= "000000";
				when "000010000001100000" => data <= "000000";
				when "000010000001100001" => data <= "000000";
				when "000010000001100010" => data <= "000000";
				when "000010000001100011" => data <= "000000";
				when "000010000001100100" => data <= "000000";
				when "000010000001100101" => data <= "000000";
				when "000010000001100110" => data <= "000000";
				when "000010000001100111" => data <= "000000";
				when "000010000001101000" => data <= "000000";
				when "000010000001101001" => data <= "000000";
				when "000010000001101010" => data <= "000000";
				when "000010000001101011" => data <= "000000";
				when "000010000001101100" => data <= "000000";
				when "000010000001101101" => data <= "000000";
				when "000010000001101110" => data <= "000000";
				when "000010000001101111" => data <= "000000";
				when "000010000001110000" => data <= "000000";
				when "000010000001110001" => data <= "000000";
				when "000010000001110010" => data <= "000000";
				when "000010000001110011" => data <= "000000";
				when "000010000001110100" => data <= "000000";
				when "000010000001110101" => data <= "000000";
				when "000010000001110110" => data <= "000000";
				when "000010000001110111" => data <= "000000";
				when "000010000001111000" => data <= "000000";
				when "000010000001111001" => data <= "000000";
				when "000010000001111010" => data <= "000000";
				when "000010000001111011" => data <= "000000";
				when "000010000001111100" => data <= "000000";
				when "000010000001111101" => data <= "000000";
				when "000010000001111110" => data <= "000000";
				when "000010000001111111" => data <= "000000";
				when "000010000010000000" => data <= "000000";
				when "000010000010000001" => data <= "000000";
				when "000010000010000010" => data <= "000000";
				when "000010000010000011" => data <= "000000";
				when "000010000010000100" => data <= "000000";
				when "000010000010000101" => data <= "000000";
				when "000010000010000110" => data <= "000000";
				when "000010000010000111" => data <= "000000";
				when "000010000010001000" => data <= "000000";
				when "000010000010001001" => data <= "000000";
				when "000010000010001010" => data <= "000000";
				when "000010000010001011" => data <= "000000";
				when "000010000010001100" => data <= "000000";
				when "000010000010001101" => data <= "000000";
				when "000010000010001110" => data <= "000000";
				when "000010000010001111" => data <= "000000";
				when "000010000010010000" => data <= "000000";
				when "000010000010010001" => data <= "000000";
				when "000010000010010010" => data <= "000000";
				when "000010000010010011" => data <= "000000";
				when "000010000010010100" => data <= "000000";
				when "000010000010010101" => data <= "000000";
				when "000010000010010110" => data <= "000000";
				when "000010000010010111" => data <= "000000";
				when "000010000010011000" => data <= "000000";
				when "000010000010011001" => data <= "000000";
				when "000010000010011010" => data <= "000000";
				when "000010000010011011" => data <= "000000";
				when "000010000010011100" => data <= "000000";
				when "000010000010011101" => data <= "000000";
				when "000010000010011110" => data <= "000000";
				when "000010000010011111" => data <= "000000";
				when "000010001000000000" => data <= "000000";
				when "000010001000000001" => data <= "000000";
				when "000010001000000010" => data <= "000000";
				when "000010001000000011" => data <= "000000";
				when "000010001000000100" => data <= "000000";
				when "000010001000000101" => data <= "000000";
				when "000010001000000110" => data <= "000000";
				when "000010001000000111" => data <= "000000";
				when "000010001000001000" => data <= "000000";
				when "000010001000001001" => data <= "000000";
				when "000010001000001010" => data <= "000000";
				when "000010001000001011" => data <= "000000";
				when "000010001000001100" => data <= "000000";
				when "000010001000001101" => data <= "000000";
				when "000010001000001110" => data <= "000000";
				when "000010001000001111" => data <= "000000";
				when "000010001000010000" => data <= "000000";
				when "000010001000010001" => data <= "000000";
				when "000010001000010010" => data <= "000000";
				when "000010001000010011" => data <= "000000";
				when "000010001000010100" => data <= "000000";
				when "000010001000010101" => data <= "000000";
				when "000010001000010110" => data <= "000000";
				when "000010001000010111" => data <= "000000";
				when "000010001000011000" => data <= "000000";
				when "000010001000011001" => data <= "000000";
				when "000010001000011010" => data <= "000000";
				when "000010001000011011" => data <= "000000";
				when "000010001000011100" => data <= "000000";
				when "000010001000011101" => data <= "000000";
				when "000010001000011110" => data <= "000000";
				when "000010001000011111" => data <= "000000";
				when "000010001000100000" => data <= "000000";
				when "000010001000100001" => data <= "000000";
				when "000010001000100010" => data <= "000000";
				when "000010001000100011" => data <= "000000";
				when "000010001000100100" => data <= "000000";
				when "000010001000100101" => data <= "000000";
				when "000010001000100110" => data <= "000000";
				when "000010001000100111" => data <= "000000";
				when "000010001000101000" => data <= "000000";
				when "000010001000101001" => data <= "000000";
				when "000010001000101010" => data <= "000000";
				when "000010001000101011" => data <= "000000";
				when "000010001000101100" => data <= "000000";
				when "000010001000101101" => data <= "000000";
				when "000010001000101110" => data <= "000000";
				when "000010001000101111" => data <= "000000";
				when "000010001000110000" => data <= "000000";
				when "000010001000110001" => data <= "000000";
				when "000010001000110010" => data <= "000000";
				when "000010001000110011" => data <= "000000";
				when "000010001000110100" => data <= "000000";
				when "000010001000110101" => data <= "000000";
				when "000010001000110110" => data <= "000000";
				when "000010001000110111" => data <= "000000";
				when "000010001000111000" => data <= "000000";
				when "000010001000111001" => data <= "000000";
				when "000010001000111010" => data <= "000000";
				when "000010001000111011" => data <= "000000";
				when "000010001000111100" => data <= "000000";
				when "000010001000111101" => data <= "000000";
				when "000010001000111110" => data <= "000000";
				when "000010001000111111" => data <= "000000";
				when "000010001001000000" => data <= "000000";
				when "000010001001000001" => data <= "000000";
				when "000010001001000010" => data <= "000000";
				when "000010001001000011" => data <= "000000";
				when "000010001001000100" => data <= "000000";
				when "000010001001000101" => data <= "000000";
				when "000010001001000110" => data <= "000000";
				when "000010001001000111" => data <= "000000";
				when "000010001001001000" => data <= "000000";
				when "000010001001001001" => data <= "000000";
				when "000010001001001010" => data <= "000000";
				when "000010001001001011" => data <= "000000";
				when "000010001001001100" => data <= "000000";
				when "000010001001001101" => data <= "000000";
				when "000010001001001110" => data <= "000000";
				when "000010001001001111" => data <= "000000";
				when "000010001001010000" => data <= "000000";
				when "000010001001010001" => data <= "000000";
				when "000010001001010010" => data <= "000000";
				when "000010001001010011" => data <= "000000";
				when "000010001001010100" => data <= "000000";
				when "000010001001010101" => data <= "000000";
				when "000010001001010110" => data <= "000000";
				when "000010001001010111" => data <= "000000";
				when "000010001001011000" => data <= "000000";
				when "000010001001011001" => data <= "000000";
				when "000010001001011010" => data <= "000000";
				when "000010001001011011" => data <= "000000";
				when "000010001001011100" => data <= "000000";
				when "000010001001011101" => data <= "000000";
				when "000010001001011110" => data <= "000000";
				when "000010001001011111" => data <= "000000";
				when "000010001001100000" => data <= "000000";
				when "000010001001100001" => data <= "000000";
				when "000010001001100010" => data <= "000000";
				when "000010001001100011" => data <= "000000";
				when "000010001001100100" => data <= "000000";
				when "000010001001100101" => data <= "000000";
				when "000010001001100110" => data <= "000000";
				when "000010001001100111" => data <= "000000";
				when "000010001001101000" => data <= "000000";
				when "000010001001101001" => data <= "000000";
				when "000010001001101010" => data <= "000000";
				when "000010001001101011" => data <= "000000";
				when "000010001001101100" => data <= "000000";
				when "000010001001101101" => data <= "000000";
				when "000010001001101110" => data <= "000000";
				when "000010001001101111" => data <= "000000";
				when "000010001001110000" => data <= "000000";
				when "000010001001110001" => data <= "000000";
				when "000010001001110010" => data <= "000000";
				when "000010001001110011" => data <= "000000";
				when "000010001001110100" => data <= "000000";
				when "000010001001110101" => data <= "000000";
				when "000010001001110110" => data <= "000000";
				when "000010001001110111" => data <= "000000";
				when "000010001001111000" => data <= "000000";
				when "000010001001111001" => data <= "000000";
				when "000010001001111010" => data <= "000000";
				when "000010001001111011" => data <= "000000";
				when "000010001001111100" => data <= "000000";
				when "000010001001111101" => data <= "000000";
				when "000010001001111110" => data <= "000000";
				when "000010001001111111" => data <= "000000";
				when "000010001010000000" => data <= "000000";
				when "000010001010000001" => data <= "000000";
				when "000010001010000010" => data <= "000000";
				when "000010001010000011" => data <= "000000";
				when "000010001010000100" => data <= "000000";
				when "000010001010000101" => data <= "000000";
				when "000010001010000110" => data <= "000000";
				when "000010001010000111" => data <= "000000";
				when "000010001010001000" => data <= "000000";
				when "000010001010001001" => data <= "000000";
				when "000010001010001010" => data <= "000000";
				when "000010001010001011" => data <= "000000";
				when "000010001010001100" => data <= "000000";
				when "000010001010001101" => data <= "000000";
				when "000010001010001110" => data <= "000000";
				when "000010001010001111" => data <= "000000";
				when "000010001010010000" => data <= "000000";
				when "000010001010010001" => data <= "000000";
				when "000010001010010010" => data <= "000000";
				when "000010001010010011" => data <= "000000";
				when "000010001010010100" => data <= "000000";
				when "000010001010010101" => data <= "000000";
				when "000010001010010110" => data <= "000000";
				when "000010001010010111" => data <= "000000";
				when "000010001010011000" => data <= "000000";
				when "000010001010011001" => data <= "000000";
				when "000010001010011010" => data <= "000000";
				when "000010001010011011" => data <= "000000";
				when "000010001010011100" => data <= "000000";
				when "000010001010011101" => data <= "000000";
				when "000010001010011110" => data <= "000000";
				when "000010001010011111" => data <= "000000";
				when "000010010000000000" => data <= "000000";
				when "000010010000000001" => data <= "000000";
				when "000010010000000010" => data <= "000000";
				when "000010010000000011" => data <= "000000";
				when "000010010000000100" => data <= "000000";
				when "000010010000000101" => data <= "000000";
				when "000010010000000110" => data <= "000000";
				when "000010010000000111" => data <= "000000";
				when "000010010000001000" => data <= "000000";
				when "000010010000001001" => data <= "000000";
				when "000010010000001010" => data <= "000000";
				when "000010010000001011" => data <= "000000";
				when "000010010000001100" => data <= "000000";
				when "000010010000001101" => data <= "000000";
				when "000010010000001110" => data <= "000000";
				when "000010010000001111" => data <= "000000";
				when "000010010000010000" => data <= "000000";
				when "000010010000010001" => data <= "000000";
				when "000010010000010010" => data <= "000000";
				when "000010010000010011" => data <= "000000";
				when "000010010000010100" => data <= "000000";
				when "000010010000010101" => data <= "000000";
				when "000010010000010110" => data <= "000000";
				when "000010010000010111" => data <= "000000";
				when "000010010000011000" => data <= "000000";
				when "000010010000011001" => data <= "000000";
				when "000010010000011010" => data <= "000000";
				when "000010010000011011" => data <= "000000";
				when "000010010000011100" => data <= "000000";
				when "000010010000011101" => data <= "000000";
				when "000010010000011110" => data <= "000000";
				when "000010010000011111" => data <= "000000";
				when "000010010000100000" => data <= "000000";
				when "000010010000100001" => data <= "000000";
				when "000010010000100010" => data <= "000000";
				when "000010010000100011" => data <= "000000";
				when "000010010000100100" => data <= "000000";
				when "000010010000100101" => data <= "000000";
				when "000010010000100110" => data <= "000000";
				when "000010010000100111" => data <= "000000";
				when "000010010000101000" => data <= "000000";
				when "000010010000101001" => data <= "000000";
				when "000010010000101010" => data <= "000000";
				when "000010010000101011" => data <= "000000";
				when "000010010000101100" => data <= "000000";
				when "000010010000101101" => data <= "000000";
				when "000010010000101110" => data <= "000000";
				when "000010010000101111" => data <= "000000";
				when "000010010000110000" => data <= "000000";
				when "000010010000110001" => data <= "000000";
				when "000010010000110010" => data <= "000000";
				when "000010010000110011" => data <= "000000";
				when "000010010000110100" => data <= "000000";
				when "000010010000110101" => data <= "000000";
				when "000010010000110110" => data <= "000000";
				when "000010010000110111" => data <= "000000";
				when "000010010000111000" => data <= "000000";
				when "000010010000111001" => data <= "000000";
				when "000010010000111010" => data <= "000000";
				when "000010010000111011" => data <= "000000";
				when "000010010000111100" => data <= "000000";
				when "000010010000111101" => data <= "000000";
				when "000010010000111110" => data <= "000000";
				when "000010010000111111" => data <= "000000";
				when "000010010001000000" => data <= "000000";
				when "000010010001000001" => data <= "000000";
				when "000010010001000010" => data <= "000000";
				when "000010010001000011" => data <= "000000";
				when "000010010001000100" => data <= "000000";
				when "000010010001000101" => data <= "000000";
				when "000010010001000110" => data <= "000000";
				when "000010010001000111" => data <= "000000";
				when "000010010001001000" => data <= "000000";
				when "000010010001001001" => data <= "000000";
				when "000010010001001010" => data <= "000000";
				when "000010010001001011" => data <= "000000";
				when "000010010001001100" => data <= "000000";
				when "000010010001001101" => data <= "000000";
				when "000010010001001110" => data <= "000000";
				when "000010010001001111" => data <= "000000";
				when "000010010001010000" => data <= "000000";
				when "000010010001010001" => data <= "000000";
				when "000010010001010010" => data <= "000000";
				when "000010010001010011" => data <= "000000";
				when "000010010001010100" => data <= "000000";
				when "000010010001010101" => data <= "000000";
				when "000010010001010110" => data <= "000000";
				when "000010010001010111" => data <= "000000";
				when "000010010001011000" => data <= "000000";
				when "000010010001011001" => data <= "000000";
				when "000010010001011010" => data <= "000000";
				when "000010010001011011" => data <= "000000";
				when "000010010001011100" => data <= "000000";
				when "000010010001011101" => data <= "000000";
				when "000010010001011110" => data <= "000000";
				when "000010010001011111" => data <= "000000";
				when "000010010001100000" => data <= "000000";
				when "000010010001100001" => data <= "000000";
				when "000010010001100010" => data <= "000000";
				when "000010010001100011" => data <= "000000";
				when "000010010001100100" => data <= "000000";
				when "000010010001100101" => data <= "000000";
				when "000010010001100110" => data <= "000000";
				when "000010010001100111" => data <= "000000";
				when "000010010001101000" => data <= "000000";
				when "000010010001101001" => data <= "000000";
				when "000010010001101010" => data <= "000000";
				when "000010010001101011" => data <= "000000";
				when "000010010001101100" => data <= "000000";
				when "000010010001101101" => data <= "000000";
				when "000010010001101110" => data <= "000000";
				when "000010010001101111" => data <= "000000";
				when "000010010001110000" => data <= "000000";
				when "000010010001110001" => data <= "000000";
				when "000010010001110010" => data <= "000000";
				when "000010010001110011" => data <= "000000";
				when "000010010001110100" => data <= "000000";
				when "000010010001110101" => data <= "000000";
				when "000010010001110110" => data <= "000000";
				when "000010010001110111" => data <= "000000";
				when "000010010001111000" => data <= "000000";
				when "000010010001111001" => data <= "000000";
				when "000010010001111010" => data <= "000000";
				when "000010010001111011" => data <= "000000";
				when "000010010001111100" => data <= "000000";
				when "000010010001111101" => data <= "000000";
				when "000010010001111110" => data <= "000000";
				when "000010010001111111" => data <= "000000";
				when "000010010010000000" => data <= "000000";
				when "000010010010000001" => data <= "000000";
				when "000010010010000010" => data <= "000000";
				when "000010010010000011" => data <= "000000";
				when "000010010010000100" => data <= "000000";
				when "000010010010000101" => data <= "000000";
				when "000010010010000110" => data <= "000000";
				when "000010010010000111" => data <= "000000";
				when "000010010010001000" => data <= "000000";
				when "000010010010001001" => data <= "000000";
				when "000010010010001010" => data <= "000000";
				when "000010010010001011" => data <= "000000";
				when "000010010010001100" => data <= "000000";
				when "000010010010001101" => data <= "000000";
				when "000010010010001110" => data <= "000000";
				when "000010010010001111" => data <= "000000";
				when "000010010010010000" => data <= "000000";
				when "000010010010010001" => data <= "000000";
				when "000010010010010010" => data <= "000000";
				when "000010010010010011" => data <= "000000";
				when "000010010010010100" => data <= "000000";
				when "000010010010010101" => data <= "000000";
				when "000010010010010110" => data <= "000000";
				when "000010010010010111" => data <= "000000";
				when "000010010010011000" => data <= "000000";
				when "000010010010011001" => data <= "000000";
				when "000010010010011010" => data <= "000000";
				when "000010010010011011" => data <= "000000";
				when "000010010010011100" => data <= "000000";
				when "000010010010011101" => data <= "000000";
				when "000010010010011110" => data <= "000000";
				when "000010010010011111" => data <= "000000";
				when "000010011000000000" => data <= "000000";
				when "000010011000000001" => data <= "000000";
				when "000010011000000010" => data <= "000000";
				when "000010011000000011" => data <= "000000";
				when "000010011000000100" => data <= "000000";
				when "000010011000000101" => data <= "000000";
				when "000010011000000110" => data <= "000000";
				when "000010011000000111" => data <= "000000";
				when "000010011000001000" => data <= "000000";
				when "000010011000001001" => data <= "000000";
				when "000010011000001010" => data <= "000000";
				when "000010011000001011" => data <= "000000";
				when "000010011000001100" => data <= "000000";
				when "000010011000001101" => data <= "000000";
				when "000010011000001110" => data <= "000000";
				when "000010011000001111" => data <= "000000";
				when "000010011000010000" => data <= "000000";
				when "000010011000010001" => data <= "000000";
				when "000010011000010010" => data <= "000000";
				when "000010011000010011" => data <= "000000";
				when "000010011000010100" => data <= "000000";
				when "000010011000010101" => data <= "000000";
				when "000010011000010110" => data <= "000000";
				when "000010011000010111" => data <= "000000";
				when "000010011000011000" => data <= "000000";
				when "000010011000011001" => data <= "000000";
				when "000010011000011010" => data <= "000000";
				when "000010011000011011" => data <= "000000";
				when "000010011000011100" => data <= "000000";
				when "000010011000011101" => data <= "000000";
				when "000010011000011110" => data <= "000000";
				when "000010011000011111" => data <= "000000";
				when "000010011000100000" => data <= "000000";
				when "000010011000100001" => data <= "000000";
				when "000010011000100010" => data <= "000000";
				when "000010011000100011" => data <= "000000";
				when "000010011000100100" => data <= "000000";
				when "000010011000100101" => data <= "000000";
				when "000010011000100110" => data <= "000000";
				when "000010011000100111" => data <= "000000";
				when "000010011000101000" => data <= "000000";
				when "000010011000101001" => data <= "000000";
				when "000010011000101010" => data <= "000000";
				when "000010011000101011" => data <= "000000";
				when "000010011000101100" => data <= "000000";
				when "000010011000101101" => data <= "000000";
				when "000010011000101110" => data <= "000000";
				when "000010011000101111" => data <= "000000";
				when "000010011000110000" => data <= "000000";
				when "000010011000110001" => data <= "000000";
				when "000010011000110010" => data <= "000000";
				when "000010011000110011" => data <= "000000";
				when "000010011000110100" => data <= "000000";
				when "000010011000110101" => data <= "000000";
				when "000010011000110110" => data <= "000000";
				when "000010011000110111" => data <= "000000";
				when "000010011000111000" => data <= "000000";
				when "000010011000111001" => data <= "000000";
				when "000010011000111010" => data <= "000000";
				when "000010011000111011" => data <= "000000";
				when "000010011000111100" => data <= "000000";
				when "000010011000111101" => data <= "000000";
				when "000010011000111110" => data <= "000000";
				when "000010011000111111" => data <= "000000";
				when "000010011001000000" => data <= "000000";
				when "000010011001000001" => data <= "000000";
				when "000010011001000010" => data <= "000000";
				when "000010011001000011" => data <= "000000";
				when "000010011001000100" => data <= "000000";
				when "000010011001000101" => data <= "000000";
				when "000010011001000110" => data <= "000000";
				when "000010011001000111" => data <= "000000";
				when "000010011001001000" => data <= "000000";
				when "000010011001001001" => data <= "000000";
				when "000010011001001010" => data <= "000000";
				when "000010011001001011" => data <= "000000";
				when "000010011001001100" => data <= "000000";
				when "000010011001001101" => data <= "000000";
				when "000010011001001110" => data <= "000000";
				when "000010011001001111" => data <= "000000";
				when "000010011001010000" => data <= "000000";
				when "000010011001010001" => data <= "000000";
				when "000010011001010010" => data <= "000000";
				when "000010011001010011" => data <= "000000";
				when "000010011001010100" => data <= "000000";
				when "000010011001010101" => data <= "000000";
				when "000010011001010110" => data <= "000000";
				when "000010011001010111" => data <= "000000";
				when "000010011001011000" => data <= "000000";
				when "000010011001011001" => data <= "000000";
				when "000010011001011010" => data <= "000000";
				when "000010011001011011" => data <= "000000";
				when "000010011001011100" => data <= "000000";
				when "000010011001011101" => data <= "000000";
				when "000010011001011110" => data <= "000000";
				when "000010011001011111" => data <= "000000";
				when "000010011001100000" => data <= "000000";
				when "000010011001100001" => data <= "000000";
				when "000010011001100010" => data <= "000000";
				when "000010011001100011" => data <= "000000";
				when "000010011001100100" => data <= "000000";
				when "000010011001100101" => data <= "000000";
				when "000010011001100110" => data <= "000000";
				when "000010011001100111" => data <= "000000";
				when "000010011001101000" => data <= "000000";
				when "000010011001101001" => data <= "000000";
				when "000010011001101010" => data <= "000000";
				when "000010011001101011" => data <= "000000";
				when "000010011001101100" => data <= "000000";
				when "000010011001101101" => data <= "000000";
				when "000010011001101110" => data <= "000000";
				when "000010011001101111" => data <= "000000";
				when "000010011001110000" => data <= "000000";
				when "000010011001110001" => data <= "000000";
				when "000010011001110010" => data <= "000000";
				when "000010011001110011" => data <= "000000";
				when "000010011001110100" => data <= "000000";
				when "000010011001110101" => data <= "000000";
				when "000010011001110110" => data <= "000000";
				when "000010011001110111" => data <= "000000";
				when "000010011001111000" => data <= "000000";
				when "000010011001111001" => data <= "000000";
				when "000010011001111010" => data <= "000000";
				when "000010011001111011" => data <= "000000";
				when "000010011001111100" => data <= "000000";
				when "000010011001111101" => data <= "000000";
				when "000010011001111110" => data <= "000000";
				when "000010011001111111" => data <= "000000";
				when "000010011010000000" => data <= "000000";
				when "000010011010000001" => data <= "000000";
				when "000010011010000010" => data <= "000000";
				when "000010011010000011" => data <= "000000";
				when "000010011010000100" => data <= "000000";
				when "000010011010000101" => data <= "000000";
				when "000010011010000110" => data <= "000000";
				when "000010011010000111" => data <= "000000";
				when "000010011010001000" => data <= "000000";
				when "000010011010001001" => data <= "000000";
				when "000010011010001010" => data <= "000000";
				when "000010011010001011" => data <= "000000";
				when "000010011010001100" => data <= "000000";
				when "000010011010001101" => data <= "000000";
				when "000010011010001110" => data <= "000000";
				when "000010011010001111" => data <= "000000";
				when "000010011010010000" => data <= "000000";
				when "000010011010010001" => data <= "000000";
				when "000010011010010010" => data <= "000000";
				when "000010011010010011" => data <= "000000";
				when "000010011010010100" => data <= "000000";
				when "000010011010010101" => data <= "000000";
				when "000010011010010110" => data <= "000000";
				when "000010011010010111" => data <= "000000";
				when "000010011010011000" => data <= "000000";
				when "000010011010011001" => data <= "000000";
				when "000010011010011010" => data <= "000000";
				when "000010011010011011" => data <= "000000";
				when "000010011010011100" => data <= "000000";
				when "000010011010011101" => data <= "000000";
				when "000010011010011110" => data <= "000000";
				when "000010011010011111" => data <= "000000";
				when "000010100000000000" => data <= "000000";
				when "000010100000000001" => data <= "000000";
				when "000010100000000010" => data <= "000000";
				when "000010100000000011" => data <= "000000";
				when "000010100000000100" => data <= "000000";
				when "000010100000000101" => data <= "000000";
				when "000010100000000110" => data <= "000000";
				when "000010100000000111" => data <= "000000";
				when "000010100000001000" => data <= "000000";
				when "000010100000001001" => data <= "000000";
				when "000010100000001010" => data <= "000000";
				when "000010100000001011" => data <= "000000";
				when "000010100000001100" => data <= "000000";
				when "000010100000001101" => data <= "000000";
				when "000010100000001110" => data <= "000000";
				when "000010100000001111" => data <= "000000";
				when "000010100000010000" => data <= "000000";
				when "000010100000010001" => data <= "000000";
				when "000010100000010010" => data <= "000000";
				when "000010100000010011" => data <= "000000";
				when "000010100000010100" => data <= "000000";
				when "000010100000010101" => data <= "000000";
				when "000010100000010110" => data <= "000000";
				when "000010100000010111" => data <= "000000";
				when "000010100000011000" => data <= "000000";
				when "000010100000011001" => data <= "000000";
				when "000010100000011010" => data <= "000000";
				when "000010100000011011" => data <= "000000";
				when "000010100000011100" => data <= "000000";
				when "000010100000011101" => data <= "000000";
				when "000010100000011110" => data <= "000000";
				when "000010100000011111" => data <= "000000";
				when "000010100000100000" => data <= "000000";
				when "000010100000100001" => data <= "000000";
				when "000010100000100010" => data <= "000000";
				when "000010100000100011" => data <= "000000";
				when "000010100000100100" => data <= "000000";
				when "000010100000100101" => data <= "000000";
				when "000010100000100110" => data <= "000000";
				when "000010100000100111" => data <= "000000";
				when "000010100000101000" => data <= "000000";
				when "000010100000101001" => data <= "000000";
				when "000010100000101010" => data <= "000000";
				when "000010100000101011" => data <= "000000";
				when "000010100000101100" => data <= "000000";
				when "000010100000101101" => data <= "000000";
				when "000010100000101110" => data <= "000000";
				when "000010100000101111" => data <= "000000";
				when "000010100000110000" => data <= "000000";
				when "000010100000110001" => data <= "000000";
				when "000010100000110010" => data <= "000000";
				when "000010100000110011" => data <= "000000";
				when "000010100000110100" => data <= "000000";
				when "000010100000110101" => data <= "000000";
				when "000010100000110110" => data <= "000000";
				when "000010100000110111" => data <= "000000";
				when "000010100000111000" => data <= "000000";
				when "000010100000111001" => data <= "000000";
				when "000010100000111010" => data <= "000000";
				when "000010100000111011" => data <= "000000";
				when "000010100000111100" => data <= "000000";
				when "000010100000111101" => data <= "000000";
				when "000010100000111110" => data <= "000000";
				when "000010100000111111" => data <= "000000";
				when "000010100001000000" => data <= "000000";
				when "000010100001000001" => data <= "000000";
				when "000010100001000010" => data <= "000000";
				when "000010100001000011" => data <= "000000";
				when "000010100001000100" => data <= "000000";
				when "000010100001000101" => data <= "000000";
				when "000010100001000110" => data <= "000000";
				when "000010100001000111" => data <= "000000";
				when "000010100001001000" => data <= "000000";
				when "000010100001001001" => data <= "000000";
				when "000010100001001010" => data <= "000000";
				when "000010100001001011" => data <= "000000";
				when "000010100001001100" => data <= "000000";
				when "000010100001001101" => data <= "000000";
				when "000010100001001110" => data <= "000000";
				when "000010100001001111" => data <= "000000";
				when "000010100001010000" => data <= "000000";
				when "000010100001010001" => data <= "000000";
				when "000010100001010010" => data <= "000000";
				when "000010100001010011" => data <= "000000";
				when "000010100001010100" => data <= "000000";
				when "000010100001010101" => data <= "000000";
				when "000010100001010110" => data <= "000000";
				when "000010100001010111" => data <= "000000";
				when "000010100001011000" => data <= "000000";
				when "000010100001011001" => data <= "000000";
				when "000010100001011010" => data <= "000000";
				when "000010100001011011" => data <= "000000";
				when "000010100001011100" => data <= "000000";
				when "000010100001011101" => data <= "000000";
				when "000010100001011110" => data <= "000000";
				when "000010100001011111" => data <= "000000";
				when "000010100001100000" => data <= "000000";
				when "000010100001100001" => data <= "000000";
				when "000010100001100010" => data <= "000000";
				when "000010100001100011" => data <= "000000";
				when "000010100001100100" => data <= "000000";
				when "000010100001100101" => data <= "000000";
				when "000010100001100110" => data <= "000000";
				when "000010100001100111" => data <= "000000";
				when "000010100001101000" => data <= "000000";
				when "000010100001101001" => data <= "000000";
				when "000010100001101010" => data <= "000000";
				when "000010100001101011" => data <= "000000";
				when "000010100001101100" => data <= "000000";
				when "000010100001101101" => data <= "000000";
				when "000010100001101110" => data <= "000000";
				when "000010100001101111" => data <= "000000";
				when "000010100001110000" => data <= "000000";
				when "000010100001110001" => data <= "000000";
				when "000010100001110010" => data <= "000000";
				when "000010100001110011" => data <= "000000";
				when "000010100001110100" => data <= "000000";
				when "000010100001110101" => data <= "000000";
				when "000010100001110110" => data <= "000000";
				when "000010100001110111" => data <= "000000";
				when "000010100001111000" => data <= "000000";
				when "000010100001111001" => data <= "000000";
				when "000010100001111010" => data <= "000000";
				when "000010100001111011" => data <= "000000";
				when "000010100001111100" => data <= "000000";
				when "000010100001111101" => data <= "000000";
				when "000010100001111110" => data <= "000000";
				when "000010100001111111" => data <= "000000";
				when "000010100010000000" => data <= "000000";
				when "000010100010000001" => data <= "000000";
				when "000010100010000010" => data <= "000000";
				when "000010100010000011" => data <= "000000";
				when "000010100010000100" => data <= "000000";
				when "000010100010000101" => data <= "000000";
				when "000010100010000110" => data <= "000000";
				when "000010100010000111" => data <= "000000";
				when "000010100010001000" => data <= "000000";
				when "000010100010001001" => data <= "000000";
				when "000010100010001010" => data <= "000000";
				when "000010100010001011" => data <= "000000";
				when "000010100010001100" => data <= "000000";
				when "000010100010001101" => data <= "000000";
				when "000010100010001110" => data <= "000000";
				when "000010100010001111" => data <= "000000";
				when "000010100010010000" => data <= "000000";
				when "000010100010010001" => data <= "000000";
				when "000010100010010010" => data <= "000000";
				when "000010100010010011" => data <= "000000";
				when "000010100010010100" => data <= "000000";
				when "000010100010010101" => data <= "000000";
				when "000010100010010110" => data <= "000000";
				when "000010100010010111" => data <= "000000";
				when "000010100010011000" => data <= "000000";
				when "000010100010011001" => data <= "000000";
				when "000010100010011010" => data <= "000000";
				when "000010100010011011" => data <= "000000";
				when "000010100010011100" => data <= "000000";
				when "000010100010011101" => data <= "000000";
				when "000010100010011110" => data <= "000000";
				when "000010100010011111" => data <= "000000";
				when "000010101000000000" => data <= "000000";
				when "000010101000000001" => data <= "000000";
				when "000010101000000010" => data <= "000000";
				when "000010101000000011" => data <= "000000";
				when "000010101000000100" => data <= "000000";
				when "000010101000000101" => data <= "000000";
				when "000010101000000110" => data <= "000000";
				when "000010101000000111" => data <= "000000";
				when "000010101000001000" => data <= "000000";
				when "000010101000001001" => data <= "000000";
				when "000010101000001010" => data <= "000000";
				when "000010101000001011" => data <= "000000";
				when "000010101000001100" => data <= "000000";
				when "000010101000001101" => data <= "000000";
				when "000010101000001110" => data <= "000000";
				when "000010101000001111" => data <= "000000";
				when "000010101000010000" => data <= "000000";
				when "000010101000010001" => data <= "000000";
				when "000010101000010010" => data <= "000000";
				when "000010101000010011" => data <= "000000";
				when "000010101000010100" => data <= "000000";
				when "000010101000010101" => data <= "000000";
				when "000010101000010110" => data <= "000000";
				when "000010101000010111" => data <= "000000";
				when "000010101000011000" => data <= "000000";
				when "000010101000011001" => data <= "000000";
				when "000010101000011010" => data <= "000000";
				when "000010101000011011" => data <= "000000";
				when "000010101000011100" => data <= "000000";
				when "000010101000011101" => data <= "000000";
				when "000010101000011110" => data <= "000000";
				when "000010101000011111" => data <= "000000";
				when "000010101000100000" => data <= "000000";
				when "000010101000100001" => data <= "000000";
				when "000010101000100010" => data <= "000000";
				when "000010101000100011" => data <= "000000";
				when "000010101000100100" => data <= "000000";
				when "000010101000100101" => data <= "000000";
				when "000010101000100110" => data <= "000000";
				when "000010101000100111" => data <= "000000";
				when "000010101000101000" => data <= "000000";
				when "000010101000101001" => data <= "000000";
				when "000010101000101010" => data <= "000000";
				when "000010101000101011" => data <= "000000";
				when "000010101000101100" => data <= "000000";
				when "000010101000101101" => data <= "000000";
				when "000010101000101110" => data <= "000000";
				when "000010101000101111" => data <= "000000";
				when "000010101000110000" => data <= "000000";
				when "000010101000110001" => data <= "000000";
				when "000010101000110010" => data <= "000000";
				when "000010101000110011" => data <= "000000";
				when "000010101000110100" => data <= "000000";
				when "000010101000110101" => data <= "000000";
				when "000010101000110110" => data <= "000000";
				when "000010101000110111" => data <= "000000";
				when "000010101000111000" => data <= "000000";
				when "000010101000111001" => data <= "000000";
				when "000010101000111010" => data <= "000000";
				when "000010101000111011" => data <= "000000";
				when "000010101000111100" => data <= "000000";
				when "000010101000111101" => data <= "000000";
				when "000010101000111110" => data <= "000000";
				when "000010101000111111" => data <= "000000";
				when "000010101001000000" => data <= "000000";
				when "000010101001000001" => data <= "000000";
				when "000010101001000010" => data <= "000000";
				when "000010101001000011" => data <= "000000";
				when "000010101001000100" => data <= "000000";
				when "000010101001000101" => data <= "000000";
				when "000010101001000110" => data <= "000000";
				when "000010101001000111" => data <= "000000";
				when "000010101001001000" => data <= "000000";
				when "000010101001001001" => data <= "000000";
				when "000010101001001010" => data <= "000000";
				when "000010101001001011" => data <= "000000";
				when "000010101001001100" => data <= "000000";
				when "000010101001001101" => data <= "000000";
				when "000010101001001110" => data <= "000000";
				when "000010101001001111" => data <= "000000";
				when "000010101001010000" => data <= "000000";
				when "000010101001010001" => data <= "000000";
				when "000010101001010010" => data <= "000000";
				when "000010101001010011" => data <= "000000";
				when "000010101001010100" => data <= "000000";
				when "000010101001010101" => data <= "000000";
				when "000010101001010110" => data <= "000000";
				when "000010101001010111" => data <= "000000";
				when "000010101001011000" => data <= "000000";
				when "000010101001011001" => data <= "000000";
				when "000010101001011010" => data <= "000000";
				when "000010101001011011" => data <= "000000";
				when "000010101001011100" => data <= "000000";
				when "000010101001011101" => data <= "000000";
				when "000010101001011110" => data <= "000000";
				when "000010101001011111" => data <= "000000";
				when "000010101001100000" => data <= "000000";
				when "000010101001100001" => data <= "000000";
				when "000010101001100010" => data <= "000000";
				when "000010101001100011" => data <= "000000";
				when "000010101001100100" => data <= "000000";
				when "000010101001100101" => data <= "000000";
				when "000010101001100110" => data <= "000000";
				when "000010101001100111" => data <= "000000";
				when "000010101001101000" => data <= "000000";
				when "000010101001101001" => data <= "000000";
				when "000010101001101010" => data <= "000000";
				when "000010101001101011" => data <= "000000";
				when "000010101001101100" => data <= "000000";
				when "000010101001101101" => data <= "000000";
				when "000010101001101110" => data <= "000000";
				when "000010101001101111" => data <= "000000";
				when "000010101001110000" => data <= "000000";
				when "000010101001110001" => data <= "000000";
				when "000010101001110010" => data <= "000000";
				when "000010101001110011" => data <= "000000";
				when "000010101001110100" => data <= "000000";
				when "000010101001110101" => data <= "000000";
				when "000010101001110110" => data <= "000000";
				when "000010101001110111" => data <= "000000";
				when "000010101001111000" => data <= "000000";
				when "000010101001111001" => data <= "000000";
				when "000010101001111010" => data <= "000000";
				when "000010101001111011" => data <= "000000";
				when "000010101001111100" => data <= "000000";
				when "000010101001111101" => data <= "000000";
				when "000010101001111110" => data <= "000000";
				when "000010101001111111" => data <= "000000";
				when "000010101010000000" => data <= "000000";
				when "000010101010000001" => data <= "000000";
				when "000010101010000010" => data <= "000000";
				when "000010101010000011" => data <= "000000";
				when "000010101010000100" => data <= "000000";
				when "000010101010000101" => data <= "000000";
				when "000010101010000110" => data <= "000000";
				when "000010101010000111" => data <= "000000";
				when "000010101010001000" => data <= "000000";
				when "000010101010001001" => data <= "000000";
				when "000010101010001010" => data <= "000000";
				when "000010101010001011" => data <= "000000";
				when "000010101010001100" => data <= "000000";
				when "000010101010001101" => data <= "000000";
				when "000010101010001110" => data <= "000000";
				when "000010101010001111" => data <= "000000";
				when "000010101010010000" => data <= "000000";
				when "000010101010010001" => data <= "000000";
				when "000010101010010010" => data <= "000000";
				when "000010101010010011" => data <= "000000";
				when "000010101010010100" => data <= "000000";
				when "000010101010010101" => data <= "000000";
				when "000010101010010110" => data <= "000000";
				when "000010101010010111" => data <= "000000";
				when "000010101010011000" => data <= "000000";
				when "000010101010011001" => data <= "000000";
				when "000010101010011010" => data <= "000000";
				when "000010101010011011" => data <= "000000";
				when "000010101010011100" => data <= "000000";
				when "000010101010011101" => data <= "000000";
				when "000010101010011110" => data <= "000000";
				when "000010101010011111" => data <= "000000";
				when "000010110000000000" => data <= "000000";
				when "000010110000000001" => data <= "000000";
				when "000010110000000010" => data <= "000000";
				when "000010110000000011" => data <= "000000";
				when "000010110000000100" => data <= "000000";
				when "000010110000000101" => data <= "000000";
				when "000010110000000110" => data <= "000000";
				when "000010110000000111" => data <= "000000";
				when "000010110000001000" => data <= "000000";
				when "000010110000001001" => data <= "000000";
				when "000010110000001010" => data <= "000000";
				when "000010110000001011" => data <= "000000";
				when "000010110000001100" => data <= "000000";
				when "000010110000001101" => data <= "000000";
				when "000010110000001110" => data <= "000000";
				when "000010110000001111" => data <= "000000";
				when "000010110000010000" => data <= "000000";
				when "000010110000010001" => data <= "000000";
				when "000010110000010010" => data <= "000000";
				when "000010110000010011" => data <= "000000";
				when "000010110000010100" => data <= "000000";
				when "000010110000010101" => data <= "000000";
				when "000010110000010110" => data <= "000000";
				when "000010110000010111" => data <= "000000";
				when "000010110000011000" => data <= "000000";
				when "000010110000011001" => data <= "000000";
				when "000010110000011010" => data <= "000000";
				when "000010110000011011" => data <= "000000";
				when "000010110000011100" => data <= "000000";
				when "000010110000011101" => data <= "000000";
				when "000010110000011110" => data <= "000000";
				when "000010110000011111" => data <= "000000";
				when "000010110000100000" => data <= "000000";
				when "000010110000100001" => data <= "000000";
				when "000010110000100010" => data <= "000000";
				when "000010110000100011" => data <= "000000";
				when "000010110000100100" => data <= "000000";
				when "000010110000100101" => data <= "000000";
				when "000010110000100110" => data <= "000000";
				when "000010110000100111" => data <= "000000";
				when "000010110000101000" => data <= "000000";
				when "000010110000101001" => data <= "000000";
				when "000010110000101010" => data <= "000000";
				when "000010110000101011" => data <= "000000";
				when "000010110000101100" => data <= "000000";
				when "000010110000101101" => data <= "000000";
				when "000010110000101110" => data <= "000000";
				when "000010110000101111" => data <= "000000";
				when "000010110000110000" => data <= "000000";
				when "000010110000110001" => data <= "000000";
				when "000010110000110010" => data <= "000000";
				when "000010110000110011" => data <= "000000";
				when "000010110000110100" => data <= "000000";
				when "000010110000110101" => data <= "000000";
				when "000010110000110110" => data <= "000000";
				when "000010110000110111" => data <= "000000";
				when "000010110000111000" => data <= "000000";
				when "000010110000111001" => data <= "000000";
				when "000010110000111010" => data <= "000000";
				when "000010110000111011" => data <= "000000";
				when "000010110000111100" => data <= "000000";
				when "000010110000111101" => data <= "000000";
				when "000010110000111110" => data <= "000000";
				when "000010110000111111" => data <= "000000";
				when "000010110001000000" => data <= "000000";
				when "000010110001000001" => data <= "000000";
				when "000010110001000010" => data <= "000000";
				when "000010110001000011" => data <= "000000";
				when "000010110001000100" => data <= "000000";
				when "000010110001000101" => data <= "000000";
				when "000010110001000110" => data <= "000000";
				when "000010110001000111" => data <= "000000";
				when "000010110001001000" => data <= "000000";
				when "000010110001001001" => data <= "000000";
				when "000010110001001010" => data <= "000000";
				when "000010110001001011" => data <= "000000";
				when "000010110001001100" => data <= "000000";
				when "000010110001001101" => data <= "000000";
				when "000010110001001110" => data <= "000000";
				when "000010110001001111" => data <= "000000";
				when "000010110001010000" => data <= "000000";
				when "000010110001010001" => data <= "000000";
				when "000010110001010010" => data <= "000000";
				when "000010110001010011" => data <= "000000";
				when "000010110001010100" => data <= "000000";
				when "000010110001010101" => data <= "000000";
				when "000010110001010110" => data <= "000000";
				when "000010110001010111" => data <= "000000";
				when "000010110001011000" => data <= "000000";
				when "000010110001011001" => data <= "000000";
				when "000010110001011010" => data <= "000000";
				when "000010110001011011" => data <= "000000";
				when "000010110001011100" => data <= "000000";
				when "000010110001011101" => data <= "000000";
				when "000010110001011110" => data <= "000000";
				when "000010110001011111" => data <= "000000";
				when "000010110001100000" => data <= "000000";
				when "000010110001100001" => data <= "000000";
				when "000010110001100010" => data <= "000000";
				when "000010110001100011" => data <= "000000";
				when "000010110001100100" => data <= "000000";
				when "000010110001100101" => data <= "000000";
				when "000010110001100110" => data <= "000000";
				when "000010110001100111" => data <= "000000";
				when "000010110001101000" => data <= "000000";
				when "000010110001101001" => data <= "000000";
				when "000010110001101010" => data <= "000000";
				when "000010110001101011" => data <= "000000";
				when "000010110001101100" => data <= "000000";
				when "000010110001101101" => data <= "000000";
				when "000010110001101110" => data <= "000000";
				when "000010110001101111" => data <= "000000";
				when "000010110001110000" => data <= "000000";
				when "000010110001110001" => data <= "000000";
				when "000010110001110010" => data <= "000000";
				when "000010110001110011" => data <= "000000";
				when "000010110001110100" => data <= "000000";
				when "000010110001110101" => data <= "000000";
				when "000010110001110110" => data <= "000000";
				when "000010110001110111" => data <= "000000";
				when "000010110001111000" => data <= "000000";
				when "000010110001111001" => data <= "000000";
				when "000010110001111010" => data <= "000000";
				when "000010110001111011" => data <= "000000";
				when "000010110001111100" => data <= "000000";
				when "000010110001111101" => data <= "000000";
				when "000010110001111110" => data <= "000000";
				when "000010110001111111" => data <= "000000";
				when "000010110010000000" => data <= "000000";
				when "000010110010000001" => data <= "000000";
				when "000010110010000010" => data <= "000000";
				when "000010110010000011" => data <= "000000";
				when "000010110010000100" => data <= "000000";
				when "000010110010000101" => data <= "000000";
				when "000010110010000110" => data <= "000000";
				when "000010110010000111" => data <= "000000";
				when "000010110010001000" => data <= "000000";
				when "000010110010001001" => data <= "000000";
				when "000010110010001010" => data <= "000000";
				when "000010110010001011" => data <= "000000";
				when "000010110010001100" => data <= "000000";
				when "000010110010001101" => data <= "000000";
				when "000010110010001110" => data <= "000000";
				when "000010110010001111" => data <= "000000";
				when "000010110010010000" => data <= "000000";
				when "000010110010010001" => data <= "000000";
				when "000010110010010010" => data <= "000000";
				when "000010110010010011" => data <= "000000";
				when "000010110010010100" => data <= "000000";
				when "000010110010010101" => data <= "000000";
				when "000010110010010110" => data <= "000000";
				when "000010110010010111" => data <= "000000";
				when "000010110010011000" => data <= "000000";
				when "000010110010011001" => data <= "000000";
				when "000010110010011010" => data <= "000000";
				when "000010110010011011" => data <= "000000";
				when "000010110010011100" => data <= "000000";
				when "000010110010011101" => data <= "000000";
				when "000010110010011110" => data <= "000000";
				when "000010110010011111" => data <= "000000";
				when "000010111000000000" => data <= "000000";
				when "000010111000000001" => data <= "000000";
				when "000010111000000010" => data <= "000000";
				when "000010111000000011" => data <= "000000";
				when "000010111000000100" => data <= "000000";
				when "000010111000000101" => data <= "000000";
				when "000010111000000110" => data <= "000000";
				when "000010111000000111" => data <= "000000";
				when "000010111000001000" => data <= "000000";
				when "000010111000001001" => data <= "000000";
				when "000010111000001010" => data <= "000000";
				when "000010111000001011" => data <= "000000";
				when "000010111000001100" => data <= "000000";
				when "000010111000001101" => data <= "000000";
				when "000010111000001110" => data <= "000000";
				when "000010111000001111" => data <= "000000";
				when "000010111000010000" => data <= "000000";
				when "000010111000010001" => data <= "000000";
				when "000010111000010010" => data <= "000000";
				when "000010111000010011" => data <= "000000";
				when "000010111000010100" => data <= "000000";
				when "000010111000010101" => data <= "000000";
				when "000010111000010110" => data <= "000000";
				when "000010111000010111" => data <= "000000";
				when "000010111000011000" => data <= "000000";
				when "000010111000011001" => data <= "000000";
				when "000010111000011010" => data <= "000000";
				when "000010111000011011" => data <= "000000";
				when "000010111000011100" => data <= "000000";
				when "000010111000011101" => data <= "000000";
				when "000010111000011110" => data <= "000000";
				when "000010111000011111" => data <= "000000";
				when "000010111000100000" => data <= "000000";
				when "000010111000100001" => data <= "000000";
				when "000010111000100010" => data <= "000000";
				when "000010111000100011" => data <= "000000";
				when "000010111000100100" => data <= "000000";
				when "000010111000100101" => data <= "000000";
				when "000010111000100110" => data <= "000000";
				when "000010111000100111" => data <= "000000";
				when "000010111000101000" => data <= "000000";
				when "000010111000101001" => data <= "000000";
				when "000010111000101010" => data <= "000000";
				when "000010111000101011" => data <= "000000";
				when "000010111000101100" => data <= "000000";
				when "000010111000101101" => data <= "000000";
				when "000010111000101110" => data <= "000000";
				when "000010111000101111" => data <= "000000";
				when "000010111000110000" => data <= "000000";
				when "000010111000110001" => data <= "000000";
				when "000010111000110010" => data <= "000000";
				when "000010111000110011" => data <= "000000";
				when "000010111000110100" => data <= "000000";
				when "000010111000110101" => data <= "000000";
				when "000010111000110110" => data <= "000000";
				when "000010111000110111" => data <= "000000";
				when "000010111000111000" => data <= "000000";
				when "000010111000111001" => data <= "000000";
				when "000010111000111010" => data <= "000000";
				when "000010111000111011" => data <= "000000";
				when "000010111000111100" => data <= "000000";
				when "000010111000111101" => data <= "000000";
				when "000010111000111110" => data <= "000000";
				when "000010111000111111" => data <= "000000";
				when "000010111001000000" => data <= "000000";
				when "000010111001000001" => data <= "000000";
				when "000010111001000010" => data <= "000000";
				when "000010111001000011" => data <= "000000";
				when "000010111001000100" => data <= "000000";
				when "000010111001000101" => data <= "000000";
				when "000010111001000110" => data <= "000000";
				when "000010111001000111" => data <= "000000";
				when "000010111001001000" => data <= "000000";
				when "000010111001001001" => data <= "000000";
				when "000010111001001010" => data <= "000000";
				when "000010111001001011" => data <= "000000";
				when "000010111001001100" => data <= "000000";
				when "000010111001001101" => data <= "000000";
				when "000010111001001110" => data <= "000000";
				when "000010111001001111" => data <= "000000";
				when "000010111001010000" => data <= "000000";
				when "000010111001010001" => data <= "000000";
				when "000010111001010010" => data <= "000000";
				when "000010111001010011" => data <= "000000";
				when "000010111001010100" => data <= "000000";
				when "000010111001010101" => data <= "000000";
				when "000010111001010110" => data <= "000000";
				when "000010111001010111" => data <= "000000";
				when "000010111001011000" => data <= "000000";
				when "000010111001011001" => data <= "000000";
				when "000010111001011010" => data <= "000000";
				when "000010111001011011" => data <= "000000";
				when "000010111001011100" => data <= "000000";
				when "000010111001011101" => data <= "000000";
				when "000010111001011110" => data <= "000000";
				when "000010111001011111" => data <= "000000";
				when "000010111001100000" => data <= "000000";
				when "000010111001100001" => data <= "000000";
				when "000010111001100010" => data <= "000000";
				when "000010111001100011" => data <= "000000";
				when "000010111001100100" => data <= "000000";
				when "000010111001100101" => data <= "000000";
				when "000010111001100110" => data <= "000000";
				when "000010111001100111" => data <= "000000";
				when "000010111001101000" => data <= "000000";
				when "000010111001101001" => data <= "000000";
				when "000010111001101010" => data <= "000000";
				when "000010111001101011" => data <= "000000";
				when "000010111001101100" => data <= "000000";
				when "000010111001101101" => data <= "000000";
				when "000010111001101110" => data <= "000000";
				when "000010111001101111" => data <= "000000";
				when "000010111001110000" => data <= "000000";
				when "000010111001110001" => data <= "000000";
				when "000010111001110010" => data <= "000000";
				when "000010111001110011" => data <= "000000";
				when "000010111001110100" => data <= "000000";
				when "000010111001110101" => data <= "000000";
				when "000010111001110110" => data <= "000000";
				when "000010111001110111" => data <= "000000";
				when "000010111001111000" => data <= "000000";
				when "000010111001111001" => data <= "000000";
				when "000010111001111010" => data <= "000000";
				when "000010111001111011" => data <= "000000";
				when "000010111001111100" => data <= "000000";
				when "000010111001111101" => data <= "000000";
				when "000010111001111110" => data <= "000000";
				when "000010111001111111" => data <= "000000";
				when "000010111010000000" => data <= "000000";
				when "000010111010000001" => data <= "000000";
				when "000010111010000010" => data <= "000000";
				when "000010111010000011" => data <= "000000";
				when "000010111010000100" => data <= "000000";
				when "000010111010000101" => data <= "000000";
				when "000010111010000110" => data <= "000000";
				when "000010111010000111" => data <= "000000";
				when "000010111010001000" => data <= "000000";
				when "000010111010001001" => data <= "000000";
				when "000010111010001010" => data <= "000000";
				when "000010111010001011" => data <= "000000";
				when "000010111010001100" => data <= "000000";
				when "000010111010001101" => data <= "000000";
				when "000010111010001110" => data <= "000000";
				when "000010111010001111" => data <= "000000";
				when "000010111010010000" => data <= "000000";
				when "000010111010010001" => data <= "000000";
				when "000010111010010010" => data <= "000000";
				when "000010111010010011" => data <= "000000";
				when "000010111010010100" => data <= "000000";
				when "000010111010010101" => data <= "000000";
				when "000010111010010110" => data <= "000000";
				when "000010111010010111" => data <= "000000";
				when "000010111010011000" => data <= "000000";
				when "000010111010011001" => data <= "000000";
				when "000010111010011010" => data <= "000000";
				when "000010111010011011" => data <= "000000";
				when "000010111010011100" => data <= "000000";
				when "000010111010011101" => data <= "000000";
				when "000010111010011110" => data <= "000000";
				when "000010111010011111" => data <= "000000";
				when "000011000000000000" => data <= "000000";
				when "000011000000000001" => data <= "000000";
				when "000011000000000010" => data <= "000000";
				when "000011000000000011" => data <= "000000";
				when "000011000000000100" => data <= "000000";
				when "000011000000000101" => data <= "000000";
				when "000011000000000110" => data <= "000000";
				when "000011000000000111" => data <= "000000";
				when "000011000000001000" => data <= "000000";
				when "000011000000001001" => data <= "000000";
				when "000011000000001010" => data <= "000000";
				when "000011000000001011" => data <= "000000";
				when "000011000000001100" => data <= "000000";
				when "000011000000001101" => data <= "000000";
				when "000011000000001110" => data <= "000000";
				when "000011000000001111" => data <= "000000";
				when "000011000000010000" => data <= "000000";
				when "000011000000010001" => data <= "000000";
				when "000011000000010010" => data <= "000000";
				when "000011000000010011" => data <= "000000";
				when "000011000000010100" => data <= "000000";
				when "000011000000010101" => data <= "000000";
				when "000011000000010110" => data <= "000000";
				when "000011000000010111" => data <= "000000";
				when "000011000000011000" => data <= "000000";
				when "000011000000011001" => data <= "000000";
				when "000011000000011010" => data <= "000000";
				when "000011000000011011" => data <= "000000";
				when "000011000000011100" => data <= "000000";
				when "000011000000011101" => data <= "000000";
				when "000011000000011110" => data <= "000000";
				when "000011000000011111" => data <= "000000";
				when "000011000000100000" => data <= "000000";
				when "000011000000100001" => data <= "000000";
				when "000011000000100010" => data <= "000000";
				when "000011000000100011" => data <= "000000";
				when "000011000000100100" => data <= "000000";
				when "000011000000100101" => data <= "000000";
				when "000011000000100110" => data <= "000000";
				when "000011000000100111" => data <= "000000";
				when "000011000000101000" => data <= "000000";
				when "000011000000101001" => data <= "000000";
				when "000011000000101010" => data <= "000000";
				when "000011000000101011" => data <= "000000";
				when "000011000000101100" => data <= "000000";
				when "000011000000101101" => data <= "000000";
				when "000011000000101110" => data <= "000000";
				when "000011000000101111" => data <= "000000";
				when "000011000000110000" => data <= "000000";
				when "000011000000110001" => data <= "000000";
				when "000011000000110010" => data <= "000000";
				when "000011000000110011" => data <= "000000";
				when "000011000000110100" => data <= "000000";
				when "000011000000110101" => data <= "000000";
				when "000011000000110110" => data <= "000000";
				when "000011000000110111" => data <= "000000";
				when "000011000000111000" => data <= "000000";
				when "000011000000111001" => data <= "000000";
				when "000011000000111010" => data <= "000000";
				when "000011000000111011" => data <= "000000";
				when "000011000000111100" => data <= "000000";
				when "000011000000111101" => data <= "000000";
				when "000011000000111110" => data <= "000000";
				when "000011000000111111" => data <= "000000";
				when "000011000001000000" => data <= "000000";
				when "000011000001000001" => data <= "000000";
				when "000011000001000010" => data <= "000000";
				when "000011000001000011" => data <= "000000";
				when "000011000001000100" => data <= "000000";
				when "000011000001000101" => data <= "000000";
				when "000011000001000110" => data <= "000000";
				when "000011000001000111" => data <= "000000";
				when "000011000001001000" => data <= "000000";
				when "000011000001001001" => data <= "000000";
				when "000011000001001010" => data <= "000000";
				when "000011000001001011" => data <= "000000";
				when "000011000001001100" => data <= "000000";
				when "000011000001001101" => data <= "000000";
				when "000011000001001110" => data <= "000000";
				when "000011000001001111" => data <= "000000";
				when "000011000001010000" => data <= "000000";
				when "000011000001010001" => data <= "000000";
				when "000011000001010010" => data <= "000000";
				when "000011000001010011" => data <= "000000";
				when "000011000001010100" => data <= "000000";
				when "000011000001010101" => data <= "000000";
				when "000011000001010110" => data <= "000000";
				when "000011000001010111" => data <= "000000";
				when "000011000001011000" => data <= "000000";
				when "000011000001011001" => data <= "000000";
				when "000011000001011010" => data <= "000000";
				when "000011000001011011" => data <= "000000";
				when "000011000001011100" => data <= "000000";
				when "000011000001011101" => data <= "000000";
				when "000011000001011110" => data <= "000000";
				when "000011000001011111" => data <= "000000";
				when "000011000001100000" => data <= "000000";
				when "000011000001100001" => data <= "000000";
				when "000011000001100010" => data <= "000000";
				when "000011000001100011" => data <= "000000";
				when "000011000001100100" => data <= "000000";
				when "000011000001100101" => data <= "000000";
				when "000011000001100110" => data <= "000000";
				when "000011000001100111" => data <= "000000";
				when "000011000001101000" => data <= "000000";
				when "000011000001101001" => data <= "000000";
				when "000011000001101010" => data <= "000000";
				when "000011000001101011" => data <= "000000";
				when "000011000001101100" => data <= "000000";
				when "000011000001101101" => data <= "000000";
				when "000011000001101110" => data <= "000000";
				when "000011000001101111" => data <= "000000";
				when "000011000001110000" => data <= "000000";
				when "000011000001110001" => data <= "000000";
				when "000011000001110010" => data <= "000000";
				when "000011000001110011" => data <= "000000";
				when "000011000001110100" => data <= "000000";
				when "000011000001110101" => data <= "000000";
				when "000011000001110110" => data <= "000000";
				when "000011000001110111" => data <= "000000";
				when "000011000001111000" => data <= "000000";
				when "000011000001111001" => data <= "000000";
				when "000011000001111010" => data <= "000000";
				when "000011000001111011" => data <= "000000";
				when "000011000001111100" => data <= "000000";
				when "000011000001111101" => data <= "000000";
				when "000011000001111110" => data <= "000000";
				when "000011000001111111" => data <= "000000";
				when "000011000010000000" => data <= "000000";
				when "000011000010000001" => data <= "000000";
				when "000011000010000010" => data <= "000000";
				when "000011000010000011" => data <= "000000";
				when "000011000010000100" => data <= "000000";
				when "000011000010000101" => data <= "000000";
				when "000011000010000110" => data <= "000000";
				when "000011000010000111" => data <= "000000";
				when "000011000010001000" => data <= "000000";
				when "000011000010001001" => data <= "000000";
				when "000011000010001010" => data <= "000000";
				when "000011000010001011" => data <= "000000";
				when "000011000010001100" => data <= "000000";
				when "000011000010001101" => data <= "000000";
				when "000011000010001110" => data <= "000000";
				when "000011000010001111" => data <= "000000";
				when "000011000010010000" => data <= "000000";
				when "000011000010010001" => data <= "000000";
				when "000011000010010010" => data <= "000000";
				when "000011000010010011" => data <= "000000";
				when "000011000010010100" => data <= "000000";
				when "000011000010010101" => data <= "000000";
				when "000011000010010110" => data <= "000000";
				when "000011000010010111" => data <= "000000";
				when "000011000010011000" => data <= "000000";
				when "000011000010011001" => data <= "000000";
				when "000011000010011010" => data <= "000000";
				when "000011000010011011" => data <= "000000";
				when "000011000010011100" => data <= "000000";
				when "000011000010011101" => data <= "000000";
				when "000011000010011110" => data <= "000000";
				when "000011000010011111" => data <= "000000";
				when "000011001000000000" => data <= "000000";
				when "000011001000000001" => data <= "000000";
				when "000011001000000010" => data <= "000000";
				when "000011001000000011" => data <= "000000";
				when "000011001000000100" => data <= "000000";
				when "000011001000000101" => data <= "000000";
				when "000011001000000110" => data <= "000000";
				when "000011001000000111" => data <= "000000";
				when "000011001000001000" => data <= "000000";
				when "000011001000001001" => data <= "000000";
				when "000011001000001010" => data <= "000000";
				when "000011001000001011" => data <= "000000";
				when "000011001000001100" => data <= "000000";
				when "000011001000001101" => data <= "000000";
				when "000011001000001110" => data <= "000000";
				when "000011001000001111" => data <= "000000";
				when "000011001000010000" => data <= "000000";
				when "000011001000010001" => data <= "000000";
				when "000011001000010010" => data <= "000000";
				when "000011001000010011" => data <= "000000";
				when "000011001000010100" => data <= "000000";
				when "000011001000010101" => data <= "000000";
				when "000011001000010110" => data <= "000000";
				when "000011001000010111" => data <= "000000";
				when "000011001000011000" => data <= "000000";
				when "000011001000011001" => data <= "000000";
				when "000011001000011010" => data <= "000000";
				when "000011001000011011" => data <= "000000";
				when "000011001000011100" => data <= "000000";
				when "000011001000011101" => data <= "000000";
				when "000011001000011110" => data <= "000000";
				when "000011001000011111" => data <= "000000";
				when "000011001000100000" => data <= "000000";
				when "000011001000100001" => data <= "000000";
				when "000011001000100010" => data <= "000000";
				when "000011001000100011" => data <= "000000";
				when "000011001000100100" => data <= "000000";
				when "000011001000100101" => data <= "000000";
				when "000011001000100110" => data <= "000000";
				when "000011001000100111" => data <= "000000";
				when "000011001000101000" => data <= "000000";
				when "000011001000101001" => data <= "000000";
				when "000011001000101010" => data <= "000000";
				when "000011001000101011" => data <= "000000";
				when "000011001000101100" => data <= "000000";
				when "000011001000101101" => data <= "000000";
				when "000011001000101110" => data <= "000000";
				when "000011001000101111" => data <= "000000";
				when "000011001000110000" => data <= "000000";
				when "000011001000110001" => data <= "000000";
				when "000011001000110010" => data <= "000000";
				when "000011001000110011" => data <= "000000";
				when "000011001000110100" => data <= "000000";
				when "000011001000110101" => data <= "000000";
				when "000011001000110110" => data <= "000000";
				when "000011001000110111" => data <= "000000";
				when "000011001000111000" => data <= "000000";
				when "000011001000111001" => data <= "000000";
				when "000011001000111010" => data <= "000000";
				when "000011001000111011" => data <= "000000";
				when "000011001000111100" => data <= "000000";
				when "000011001000111101" => data <= "000000";
				when "000011001000111110" => data <= "000000";
				when "000011001000111111" => data <= "000000";
				when "000011001001000000" => data <= "000000";
				when "000011001001000001" => data <= "000000";
				when "000011001001000010" => data <= "000000";
				when "000011001001000011" => data <= "000000";
				when "000011001001000100" => data <= "000000";
				when "000011001001000101" => data <= "000000";
				when "000011001001000110" => data <= "000000";
				when "000011001001000111" => data <= "000000";
				when "000011001001001000" => data <= "000000";
				when "000011001001001001" => data <= "000000";
				when "000011001001001010" => data <= "000000";
				when "000011001001001011" => data <= "000000";
				when "000011001001001100" => data <= "000000";
				when "000011001001001101" => data <= "000000";
				when "000011001001001110" => data <= "000000";
				when "000011001001001111" => data <= "000000";
				when "000011001001010000" => data <= "000000";
				when "000011001001010001" => data <= "000000";
				when "000011001001010010" => data <= "000000";
				when "000011001001010011" => data <= "000000";
				when "000011001001010100" => data <= "000000";
				when "000011001001010101" => data <= "000000";
				when "000011001001010110" => data <= "000000";
				when "000011001001010111" => data <= "000000";
				when "000011001001011000" => data <= "000000";
				when "000011001001011001" => data <= "000000";
				when "000011001001011010" => data <= "000000";
				when "000011001001011011" => data <= "000000";
				when "000011001001011100" => data <= "000000";
				when "000011001001011101" => data <= "000000";
				when "000011001001011110" => data <= "000000";
				when "000011001001011111" => data <= "000000";
				when "000011001001100000" => data <= "000000";
				when "000011001001100001" => data <= "000000";
				when "000011001001100010" => data <= "000000";
				when "000011001001100011" => data <= "000000";
				when "000011001001100100" => data <= "000000";
				when "000011001001100101" => data <= "000000";
				when "000011001001100110" => data <= "000000";
				when "000011001001100111" => data <= "000000";
				when "000011001001101000" => data <= "000000";
				when "000011001001101001" => data <= "000000";
				when "000011001001101010" => data <= "000000";
				when "000011001001101011" => data <= "000000";
				when "000011001001101100" => data <= "000000";
				when "000011001001101101" => data <= "000000";
				when "000011001001101110" => data <= "000000";
				when "000011001001101111" => data <= "000000";
				when "000011001001110000" => data <= "000000";
				when "000011001001110001" => data <= "000000";
				when "000011001001110010" => data <= "000000";
				when "000011001001110011" => data <= "000000";
				when "000011001001110100" => data <= "000000";
				when "000011001001110101" => data <= "000000";
				when "000011001001110110" => data <= "000000";
				when "000011001001110111" => data <= "000000";
				when "000011001001111000" => data <= "000000";
				when "000011001001111001" => data <= "000000";
				when "000011001001111010" => data <= "000000";
				when "000011001001111011" => data <= "000000";
				when "000011001001111100" => data <= "000000";
				when "000011001001111101" => data <= "000000";
				when "000011001001111110" => data <= "000000";
				when "000011001001111111" => data <= "000000";
				when "000011001010000000" => data <= "000000";
				when "000011001010000001" => data <= "000000";
				when "000011001010000010" => data <= "000000";
				when "000011001010000011" => data <= "000000";
				when "000011001010000100" => data <= "000000";
				when "000011001010000101" => data <= "000000";
				when "000011001010000110" => data <= "000000";
				when "000011001010000111" => data <= "000000";
				when "000011001010001000" => data <= "000000";
				when "000011001010001001" => data <= "000000";
				when "000011001010001010" => data <= "000000";
				when "000011001010001011" => data <= "000000";
				when "000011001010001100" => data <= "000000";
				when "000011001010001101" => data <= "000000";
				when "000011001010001110" => data <= "000000";
				when "000011001010001111" => data <= "000000";
				when "000011001010010000" => data <= "000000";
				when "000011001010010001" => data <= "000000";
				when "000011001010010010" => data <= "000000";
				when "000011001010010011" => data <= "000000";
				when "000011001010010100" => data <= "000000";
				when "000011001010010101" => data <= "000000";
				when "000011001010010110" => data <= "000000";
				when "000011001010010111" => data <= "000000";
				when "000011001010011000" => data <= "000000";
				when "000011001010011001" => data <= "000000";
				when "000011001010011010" => data <= "000000";
				when "000011001010011011" => data <= "000000";
				when "000011001010011100" => data <= "000000";
				when "000011001010011101" => data <= "000000";
				when "000011001010011110" => data <= "000000";
				when "000011001010011111" => data <= "000000";
				when "000011010000000000" => data <= "000000";
				when "000011010000000001" => data <= "000000";
				when "000011010000000010" => data <= "000000";
				when "000011010000000011" => data <= "000000";
				when "000011010000000100" => data <= "000000";
				when "000011010000000101" => data <= "000000";
				when "000011010000000110" => data <= "000000";
				when "000011010000000111" => data <= "000000";
				when "000011010000001000" => data <= "000000";
				when "000011010000001001" => data <= "000000";
				when "000011010000001010" => data <= "000000";
				when "000011010000001011" => data <= "000000";
				when "000011010000001100" => data <= "000000";
				when "000011010000001101" => data <= "000000";
				when "000011010000001110" => data <= "000000";
				when "000011010000001111" => data <= "000000";
				when "000011010000010000" => data <= "000000";
				when "000011010000010001" => data <= "000000";
				when "000011010000010010" => data <= "000000";
				when "000011010000010011" => data <= "000000";
				when "000011010000010100" => data <= "000000";
				when "000011010000010101" => data <= "000000";
				when "000011010000010110" => data <= "000000";
				when "000011010000010111" => data <= "000000";
				when "000011010000011000" => data <= "000000";
				when "000011010000011001" => data <= "000000";
				when "000011010000011010" => data <= "000000";
				when "000011010000011011" => data <= "000000";
				when "000011010000011100" => data <= "000000";
				when "000011010000011101" => data <= "000000";
				when "000011010000011110" => data <= "000000";
				when "000011010000011111" => data <= "000000";
				when "000011010000100000" => data <= "000000";
				when "000011010000100001" => data <= "000000";
				when "000011010000100010" => data <= "000000";
				when "000011010000100011" => data <= "000000";
				when "000011010000100100" => data <= "000000";
				when "000011010000100101" => data <= "000000";
				when "000011010000100110" => data <= "000000";
				when "000011010000100111" => data <= "000000";
				when "000011010000101000" => data <= "000000";
				when "000011010000101001" => data <= "000000";
				when "000011010000101010" => data <= "000000";
				when "000011010000101011" => data <= "000000";
				when "000011010000101100" => data <= "000000";
				when "000011010000101101" => data <= "000000";
				when "000011010000101110" => data <= "000000";
				when "000011010000101111" => data <= "000000";
				when "000011010000110000" => data <= "000000";
				when "000011010000110001" => data <= "000000";
				when "000011010000110010" => data <= "000000";
				when "000011010000110011" => data <= "000000";
				when "000011010000110100" => data <= "000000";
				when "000011010000110101" => data <= "000000";
				when "000011010000110110" => data <= "000000";
				when "000011010000110111" => data <= "000000";
				when "000011010000111000" => data <= "000000";
				when "000011010000111001" => data <= "000000";
				when "000011010000111010" => data <= "000000";
				when "000011010000111011" => data <= "000000";
				when "000011010000111100" => data <= "000000";
				when "000011010000111101" => data <= "000000";
				when "000011010000111110" => data <= "000000";
				when "000011010000111111" => data <= "000000";
				when "000011010001000000" => data <= "000000";
				when "000011010001000001" => data <= "000000";
				when "000011010001000010" => data <= "000000";
				when "000011010001000011" => data <= "000000";
				when "000011010001000100" => data <= "000000";
				when "000011010001000101" => data <= "000000";
				when "000011010001000110" => data <= "000000";
				when "000011010001000111" => data <= "000000";
				when "000011010001001000" => data <= "000000";
				when "000011010001001001" => data <= "000000";
				when "000011010001001010" => data <= "000000";
				when "000011010001001011" => data <= "000000";
				when "000011010001001100" => data <= "000000";
				when "000011010001001101" => data <= "000000";
				when "000011010001001110" => data <= "000000";
				when "000011010001001111" => data <= "000000";
				when "000011010001010000" => data <= "000000";
				when "000011010001010001" => data <= "000000";
				when "000011010001010010" => data <= "000000";
				when "000011010001010011" => data <= "000000";
				when "000011010001010100" => data <= "000000";
				when "000011010001010101" => data <= "000000";
				when "000011010001010110" => data <= "000000";
				when "000011010001010111" => data <= "000000";
				when "000011010001011000" => data <= "000000";
				when "000011010001011001" => data <= "000000";
				when "000011010001011010" => data <= "000000";
				when "000011010001011011" => data <= "000000";
				when "000011010001011100" => data <= "000000";
				when "000011010001011101" => data <= "000000";
				when "000011010001011110" => data <= "000000";
				when "000011010001011111" => data <= "000000";
				when "000011010001100000" => data <= "000000";
				when "000011010001100001" => data <= "000000";
				when "000011010001100010" => data <= "000000";
				when "000011010001100011" => data <= "000000";
				when "000011010001100100" => data <= "000000";
				when "000011010001100101" => data <= "000000";
				when "000011010001100110" => data <= "000000";
				when "000011010001100111" => data <= "000000";
				when "000011010001101000" => data <= "000000";
				when "000011010001101001" => data <= "000000";
				when "000011010001101010" => data <= "000000";
				when "000011010001101011" => data <= "000000";
				when "000011010001101100" => data <= "000000";
				when "000011010001101101" => data <= "000000";
				when "000011010001101110" => data <= "000000";
				when "000011010001101111" => data <= "000000";
				when "000011010001110000" => data <= "000000";
				when "000011010001110001" => data <= "000000";
				when "000011010001110010" => data <= "000000";
				when "000011010001110011" => data <= "000000";
				when "000011010001110100" => data <= "000000";
				when "000011010001110101" => data <= "000000";
				when "000011010001110110" => data <= "000000";
				when "000011010001110111" => data <= "000000";
				when "000011010001111000" => data <= "000000";
				when "000011010001111001" => data <= "000000";
				when "000011010001111010" => data <= "000000";
				when "000011010001111011" => data <= "000000";
				when "000011010001111100" => data <= "000000";
				when "000011010001111101" => data <= "000000";
				when "000011010001111110" => data <= "000000";
				when "000011010001111111" => data <= "000000";
				when "000011010010000000" => data <= "000000";
				when "000011010010000001" => data <= "000000";
				when "000011010010000010" => data <= "000000";
				when "000011010010000011" => data <= "000000";
				when "000011010010000100" => data <= "000000";
				when "000011010010000101" => data <= "000000";
				when "000011010010000110" => data <= "000000";
				when "000011010010000111" => data <= "000000";
				when "000011010010001000" => data <= "000000";
				when "000011010010001001" => data <= "000000";
				when "000011010010001010" => data <= "000000";
				when "000011010010001011" => data <= "000000";
				when "000011010010001100" => data <= "000000";
				when "000011010010001101" => data <= "000000";
				when "000011010010001110" => data <= "000000";
				when "000011010010001111" => data <= "000000";
				when "000011010010010000" => data <= "000000";
				when "000011010010010001" => data <= "000000";
				when "000011010010010010" => data <= "000000";
				when "000011010010010011" => data <= "000000";
				when "000011010010010100" => data <= "000000";
				when "000011010010010101" => data <= "000000";
				when "000011010010010110" => data <= "000000";
				when "000011010010010111" => data <= "000000";
				when "000011010010011000" => data <= "000000";
				when "000011010010011001" => data <= "000000";
				when "000011010010011010" => data <= "000000";
				when "000011010010011011" => data <= "000000";
				when "000011010010011100" => data <= "000000";
				when "000011010010011101" => data <= "000000";
				when "000011010010011110" => data <= "000000";
				when "000011010010011111" => data <= "000000";
				when "000011011000000000" => data <= "000000";
				when "000011011000000001" => data <= "000000";
				when "000011011000000010" => data <= "000000";
				when "000011011000000011" => data <= "000000";
				when "000011011000000100" => data <= "000000";
				when "000011011000000101" => data <= "000000";
				when "000011011000000110" => data <= "000000";
				when "000011011000000111" => data <= "000000";
				when "000011011000001000" => data <= "000000";
				when "000011011000001001" => data <= "000000";
				when "000011011000001010" => data <= "000000";
				when "000011011000001011" => data <= "000000";
				when "000011011000001100" => data <= "000000";
				when "000011011000001101" => data <= "000000";
				when "000011011000001110" => data <= "000000";
				when "000011011000001111" => data <= "000000";
				when "000011011000010000" => data <= "000000";
				when "000011011000010001" => data <= "000000";
				when "000011011000010010" => data <= "000000";
				when "000011011000010011" => data <= "000000";
				when "000011011000010100" => data <= "000000";
				when "000011011000010101" => data <= "000000";
				when "000011011000010110" => data <= "000000";
				when "000011011000010111" => data <= "000000";
				when "000011011000011000" => data <= "000000";
				when "000011011000011001" => data <= "000000";
				when "000011011000011010" => data <= "000000";
				when "000011011000011011" => data <= "000000";
				when "000011011000011100" => data <= "000000";
				when "000011011000011101" => data <= "000000";
				when "000011011000011110" => data <= "000000";
				when "000011011000011111" => data <= "000000";
				when "000011011000100000" => data <= "000000";
				when "000011011000100001" => data <= "000000";
				when "000011011000100010" => data <= "000000";
				when "000011011000100011" => data <= "000000";
				when "000011011000100100" => data <= "000000";
				when "000011011000100101" => data <= "000000";
				when "000011011000100110" => data <= "000000";
				when "000011011000100111" => data <= "000000";
				when "000011011000101000" => data <= "000000";
				when "000011011000101001" => data <= "000000";
				when "000011011000101010" => data <= "000000";
				when "000011011000101011" => data <= "000000";
				when "000011011000101100" => data <= "000000";
				when "000011011000101101" => data <= "000000";
				when "000011011000101110" => data <= "000000";
				when "000011011000101111" => data <= "000000";
				when "000011011000110000" => data <= "000000";
				when "000011011000110001" => data <= "000000";
				when "000011011000110010" => data <= "000000";
				when "000011011000110011" => data <= "000000";
				when "000011011000110100" => data <= "000000";
				when "000011011000110101" => data <= "000000";
				when "000011011000110110" => data <= "000000";
				when "000011011000110111" => data <= "000000";
				when "000011011000111000" => data <= "000000";
				when "000011011000111001" => data <= "000000";
				when "000011011000111010" => data <= "000000";
				when "000011011000111011" => data <= "000000";
				when "000011011000111100" => data <= "000000";
				when "000011011000111101" => data <= "000000";
				when "000011011000111110" => data <= "000000";
				when "000011011000111111" => data <= "000000";
				when "000011011001000000" => data <= "000000";
				when "000011011001000001" => data <= "000000";
				when "000011011001000010" => data <= "000000";
				when "000011011001000011" => data <= "000000";
				when "000011011001000100" => data <= "000000";
				when "000011011001000101" => data <= "000000";
				when "000011011001000110" => data <= "000000";
				when "000011011001000111" => data <= "000000";
				when "000011011001001000" => data <= "000000";
				when "000011011001001001" => data <= "000000";
				when "000011011001001010" => data <= "000000";
				when "000011011001001011" => data <= "000000";
				when "000011011001001100" => data <= "000000";
				when "000011011001001101" => data <= "000000";
				when "000011011001001110" => data <= "000000";
				when "000011011001001111" => data <= "000000";
				when "000011011001010000" => data <= "000000";
				when "000011011001010001" => data <= "000000";
				when "000011011001010010" => data <= "000000";
				when "000011011001010011" => data <= "000000";
				when "000011011001010100" => data <= "000000";
				when "000011011001010101" => data <= "000000";
				when "000011011001010110" => data <= "000000";
				when "000011011001010111" => data <= "000000";
				when "000011011001011000" => data <= "000000";
				when "000011011001011001" => data <= "000000";
				when "000011011001011010" => data <= "000000";
				when "000011011001011011" => data <= "000000";
				when "000011011001011100" => data <= "000000";
				when "000011011001011101" => data <= "000000";
				when "000011011001011110" => data <= "000000";
				when "000011011001011111" => data <= "000000";
				when "000011011001100000" => data <= "000000";
				when "000011011001100001" => data <= "000000";
				when "000011011001100010" => data <= "000000";
				when "000011011001100011" => data <= "000000";
				when "000011011001100100" => data <= "000000";
				when "000011011001100101" => data <= "000000";
				when "000011011001100110" => data <= "000000";
				when "000011011001100111" => data <= "000000";
				when "000011011001101000" => data <= "000000";
				when "000011011001101001" => data <= "000000";
				when "000011011001101010" => data <= "000000";
				when "000011011001101011" => data <= "000000";
				when "000011011001101100" => data <= "000000";
				when "000011011001101101" => data <= "000000";
				when "000011011001101110" => data <= "000000";
				when "000011011001101111" => data <= "000000";
				when "000011011001110000" => data <= "000000";
				when "000011011001110001" => data <= "000000";
				when "000011011001110010" => data <= "000000";
				when "000011011001110011" => data <= "000000";
				when "000011011001110100" => data <= "000000";
				when "000011011001110101" => data <= "000000";
				when "000011011001110110" => data <= "000000";
				when "000011011001110111" => data <= "000000";
				when "000011011001111000" => data <= "000000";
				when "000011011001111001" => data <= "000000";
				when "000011011001111010" => data <= "000000";
				when "000011011001111011" => data <= "000000";
				when "000011011001111100" => data <= "000000";
				when "000011011001111101" => data <= "000000";
				when "000011011001111110" => data <= "000000";
				when "000011011001111111" => data <= "000000";
				when "000011011010000000" => data <= "000000";
				when "000011011010000001" => data <= "000000";
				when "000011011010000010" => data <= "000000";
				when "000011011010000011" => data <= "000000";
				when "000011011010000100" => data <= "000000";
				when "000011011010000101" => data <= "000000";
				when "000011011010000110" => data <= "000000";
				when "000011011010000111" => data <= "000000";
				when "000011011010001000" => data <= "000000";
				when "000011011010001001" => data <= "000000";
				when "000011011010001010" => data <= "000000";
				when "000011011010001011" => data <= "000000";
				when "000011011010001100" => data <= "000000";
				when "000011011010001101" => data <= "000000";
				when "000011011010001110" => data <= "000000";
				when "000011011010001111" => data <= "000000";
				when "000011011010010000" => data <= "000000";
				when "000011011010010001" => data <= "000000";
				when "000011011010010010" => data <= "000000";
				when "000011011010010011" => data <= "000000";
				when "000011011010010100" => data <= "000000";
				when "000011011010010101" => data <= "000000";
				when "000011011010010110" => data <= "000000";
				when "000011011010010111" => data <= "000000";
				when "000011011010011000" => data <= "000000";
				when "000011011010011001" => data <= "000000";
				when "000011011010011010" => data <= "000000";
				when "000011011010011011" => data <= "000000";
				when "000011011010011100" => data <= "000000";
				when "000011011010011101" => data <= "000000";
				when "000011011010011110" => data <= "000000";
				when "000011011010011111" => data <= "000000";
				when "000011100000000000" => data <= "000000";
				when "000011100000000001" => data <= "000000";
				when "000011100000000010" => data <= "000000";
				when "000011100000000011" => data <= "000000";
				when "000011100000000100" => data <= "000000";
				when "000011100000000101" => data <= "000000";
				when "000011100000000110" => data <= "000000";
				when "000011100000000111" => data <= "000000";
				when "000011100000001000" => data <= "000000";
				when "000011100000001001" => data <= "000000";
				when "000011100000001010" => data <= "000000";
				when "000011100000001011" => data <= "000000";
				when "000011100000001100" => data <= "000000";
				when "000011100000001101" => data <= "000000";
				when "000011100000001110" => data <= "000000";
				when "000011100000001111" => data <= "000000";
				when "000011100000010000" => data <= "000000";
				when "000011100000010001" => data <= "000000";
				when "000011100000010010" => data <= "000000";
				when "000011100000010011" => data <= "000000";
				when "000011100000010100" => data <= "000000";
				when "000011100000010101" => data <= "000000";
				when "000011100000010110" => data <= "000000";
				when "000011100000010111" => data <= "000000";
				when "000011100000011000" => data <= "000000";
				when "000011100000011001" => data <= "000000";
				when "000011100000011010" => data <= "000000";
				when "000011100000011011" => data <= "000000";
				when "000011100000011100" => data <= "000000";
				when "000011100000011101" => data <= "000000";
				when "000011100000011110" => data <= "000000";
				when "000011100000011111" => data <= "000000";
				when "000011100000100000" => data <= "000000";
				when "000011100000100001" => data <= "000000";
				when "000011100000100010" => data <= "000000";
				when "000011100000100011" => data <= "000000";
				when "000011100000100100" => data <= "000000";
				when "000011100000100101" => data <= "000000";
				when "000011100000100110" => data <= "000000";
				when "000011100000100111" => data <= "000000";
				when "000011100000101000" => data <= "000000";
				when "000011100000101001" => data <= "000000";
				when "000011100000101010" => data <= "000000";
				when "000011100000101011" => data <= "000000";
				when "000011100000101100" => data <= "000000";
				when "000011100000101101" => data <= "000000";
				when "000011100000101110" => data <= "000000";
				when "000011100000101111" => data <= "000000";
				when "000011100000110000" => data <= "000000";
				when "000011100000110001" => data <= "000000";
				when "000011100000110010" => data <= "000000";
				when "000011100000110011" => data <= "000000";
				when "000011100000110100" => data <= "000000";
				when "000011100000110101" => data <= "000000";
				when "000011100000110110" => data <= "000000";
				when "000011100000110111" => data <= "000000";
				when "000011100000111000" => data <= "000000";
				when "000011100000111001" => data <= "000000";
				when "000011100000111010" => data <= "000000";
				when "000011100000111011" => data <= "000000";
				when "000011100000111100" => data <= "000000";
				when "000011100000111101" => data <= "000000";
				when "000011100000111110" => data <= "000000";
				when "000011100000111111" => data <= "000000";
				when "000011100001000000" => data <= "000000";
				when "000011100001000001" => data <= "000000";
				when "000011100001000010" => data <= "000000";
				when "000011100001000011" => data <= "000000";
				when "000011100001000100" => data <= "000000";
				when "000011100001000101" => data <= "000000";
				when "000011100001000110" => data <= "000000";
				when "000011100001000111" => data <= "000000";
				when "000011100001001000" => data <= "000000";
				when "000011100001001001" => data <= "000000";
				when "000011100001001010" => data <= "000000";
				when "000011100001001011" => data <= "000000";
				when "000011100001001100" => data <= "000000";
				when "000011100001001101" => data <= "000000";
				when "000011100001001110" => data <= "000000";
				when "000011100001001111" => data <= "000000";
				when "000011100001010000" => data <= "000000";
				when "000011100001010001" => data <= "000000";
				when "000011100001010010" => data <= "000000";
				when "000011100001010011" => data <= "000000";
				when "000011100001010100" => data <= "000000";
				when "000011100001010101" => data <= "000000";
				when "000011100001010110" => data <= "000000";
				when "000011100001010111" => data <= "000000";
				when "000011100001011000" => data <= "000000";
				when "000011100001011001" => data <= "000000";
				when "000011100001011010" => data <= "000000";
				when "000011100001011011" => data <= "000000";
				when "000011100001011100" => data <= "000000";
				when "000011100001011101" => data <= "000000";
				when "000011100001011110" => data <= "000000";
				when "000011100001011111" => data <= "000000";
				when "000011100001100000" => data <= "000000";
				when "000011100001100001" => data <= "000000";
				when "000011100001100010" => data <= "000000";
				when "000011100001100011" => data <= "000000";
				when "000011100001100100" => data <= "000000";
				when "000011100001100101" => data <= "000000";
				when "000011100001100110" => data <= "000000";
				when "000011100001100111" => data <= "000000";
				when "000011100001101000" => data <= "000000";
				when "000011100001101001" => data <= "000000";
				when "000011100001101010" => data <= "000000";
				when "000011100001101011" => data <= "000000";
				when "000011100001101100" => data <= "000000";
				when "000011100001101101" => data <= "000000";
				when "000011100001101110" => data <= "000000";
				when "000011100001101111" => data <= "000000";
				when "000011100001110000" => data <= "000000";
				when "000011100001110001" => data <= "000000";
				when "000011100001110010" => data <= "000000";
				when "000011100001110011" => data <= "000000";
				when "000011100001110100" => data <= "000000";
				when "000011100001110101" => data <= "000000";
				when "000011100001110110" => data <= "000000";
				when "000011100001110111" => data <= "000000";
				when "000011100001111000" => data <= "000000";
				when "000011100001111001" => data <= "000000";
				when "000011100001111010" => data <= "000000";
				when "000011100001111011" => data <= "000000";
				when "000011100001111100" => data <= "000000";
				when "000011100001111101" => data <= "000000";
				when "000011100001111110" => data <= "000000";
				when "000011100001111111" => data <= "000000";
				when "000011100010000000" => data <= "000000";
				when "000011100010000001" => data <= "000000";
				when "000011100010000010" => data <= "000000";
				when "000011100010000011" => data <= "000000";
				when "000011100010000100" => data <= "000000";
				when "000011100010000101" => data <= "000000";
				when "000011100010000110" => data <= "000000";
				when "000011100010000111" => data <= "000000";
				when "000011100010001000" => data <= "000000";
				when "000011100010001001" => data <= "000000";
				when "000011100010001010" => data <= "000000";
				when "000011100010001011" => data <= "000000";
				when "000011100010001100" => data <= "000000";
				when "000011100010001101" => data <= "000000";
				when "000011100010001110" => data <= "000000";
				when "000011100010001111" => data <= "000000";
				when "000011100010010000" => data <= "000000";
				when "000011100010010001" => data <= "000000";
				when "000011100010010010" => data <= "000000";
				when "000011100010010011" => data <= "000000";
				when "000011100010010100" => data <= "000000";
				when "000011100010010101" => data <= "000000";
				when "000011100010010110" => data <= "000000";
				when "000011100010010111" => data <= "000000";
				when "000011100010011000" => data <= "000000";
				when "000011100010011001" => data <= "000000";
				when "000011100010011010" => data <= "000000";
				when "000011100010011011" => data <= "000000";
				when "000011100010011100" => data <= "000000";
				when "000011100010011101" => data <= "000000";
				when "000011100010011110" => data <= "000000";
				when "000011100010011111" => data <= "000000";
				when "000011101000000000" => data <= "000000";
				when "000011101000000001" => data <= "000000";
				when "000011101000000010" => data <= "000000";
				when "000011101000000011" => data <= "000000";
				when "000011101000000100" => data <= "000000";
				when "000011101000000101" => data <= "000000";
				when "000011101000000110" => data <= "000000";
				when "000011101000000111" => data <= "000000";
				when "000011101000001000" => data <= "000000";
				when "000011101000001001" => data <= "000000";
				when "000011101000001010" => data <= "000000";
				when "000011101000001011" => data <= "000000";
				when "000011101000001100" => data <= "000000";
				when "000011101000001101" => data <= "000000";
				when "000011101000001110" => data <= "000000";
				when "000011101000001111" => data <= "000000";
				when "000011101000010000" => data <= "000000";
				when "000011101000010001" => data <= "000000";
				when "000011101000010010" => data <= "000000";
				when "000011101000010011" => data <= "000000";
				when "000011101000010100" => data <= "000000";
				when "000011101000010101" => data <= "000000";
				when "000011101000010110" => data <= "000000";
				when "000011101000010111" => data <= "000000";
				when "000011101000011000" => data <= "000000";
				when "000011101000011001" => data <= "000000";
				when "000011101000011010" => data <= "000000";
				when "000011101000011011" => data <= "000000";
				when "000011101000011100" => data <= "000000";
				when "000011101000011101" => data <= "000000";
				when "000011101000011110" => data <= "000000";
				when "000011101000011111" => data <= "000000";
				when "000011101000100000" => data <= "000000";
				when "000011101000100001" => data <= "000000";
				when "000011101000100010" => data <= "000000";
				when "000011101000100011" => data <= "000000";
				when "000011101000100100" => data <= "000000";
				when "000011101000100101" => data <= "000000";
				when "000011101000100110" => data <= "000000";
				when "000011101000100111" => data <= "000000";
				when "000011101000101000" => data <= "000000";
				when "000011101000101001" => data <= "000000";
				when "000011101000101010" => data <= "000000";
				when "000011101000101011" => data <= "000000";
				when "000011101000101100" => data <= "000000";
				when "000011101000101101" => data <= "000000";
				when "000011101000101110" => data <= "000000";
				when "000011101000101111" => data <= "000000";
				when "000011101000110000" => data <= "000000";
				when "000011101000110001" => data <= "000000";
				when "000011101000110010" => data <= "000000";
				when "000011101000110011" => data <= "000000";
				when "000011101000110100" => data <= "000000";
				when "000011101000110101" => data <= "000000";
				when "000011101000110110" => data <= "000000";
				when "000011101000110111" => data <= "000000";
				when "000011101000111000" => data <= "000000";
				when "000011101000111001" => data <= "000000";
				when "000011101000111010" => data <= "000000";
				when "000011101000111011" => data <= "000000";
				when "000011101000111100" => data <= "000000";
				when "000011101000111101" => data <= "000000";
				when "000011101000111110" => data <= "000000";
				when "000011101000111111" => data <= "000000";
				when "000011101001000000" => data <= "000000";
				when "000011101001000001" => data <= "000000";
				when "000011101001000010" => data <= "000000";
				when "000011101001000011" => data <= "000000";
				when "000011101001000100" => data <= "000000";
				when "000011101001000101" => data <= "000000";
				when "000011101001000110" => data <= "000000";
				when "000011101001000111" => data <= "000000";
				when "000011101001001000" => data <= "000000";
				when "000011101001001001" => data <= "000000";
				when "000011101001001010" => data <= "000000";
				when "000011101001001011" => data <= "000000";
				when "000011101001001100" => data <= "000000";
				when "000011101001001101" => data <= "000000";
				when "000011101001001110" => data <= "000000";
				when "000011101001001111" => data <= "000000";
				when "000011101001010000" => data <= "000000";
				when "000011101001010001" => data <= "000000";
				when "000011101001010010" => data <= "000000";
				when "000011101001010011" => data <= "000000";
				when "000011101001010100" => data <= "000000";
				when "000011101001010101" => data <= "000000";
				when "000011101001010110" => data <= "000000";
				when "000011101001010111" => data <= "000000";
				when "000011101001011000" => data <= "000000";
				when "000011101001011001" => data <= "000000";
				when "000011101001011010" => data <= "000000";
				when "000011101001011011" => data <= "000000";
				when "000011101001011100" => data <= "000000";
				when "000011101001011101" => data <= "000000";
				when "000011101001011110" => data <= "000000";
				when "000011101001011111" => data <= "000000";
				when "000011101001100000" => data <= "000000";
				when "000011101001100001" => data <= "000000";
				when "000011101001100010" => data <= "000000";
				when "000011101001100011" => data <= "000000";
				when "000011101001100100" => data <= "000000";
				when "000011101001100101" => data <= "000000";
				when "000011101001100110" => data <= "000000";
				when "000011101001100111" => data <= "000000";
				when "000011101001101000" => data <= "000000";
				when "000011101001101001" => data <= "000000";
				when "000011101001101010" => data <= "000000";
				when "000011101001101011" => data <= "000000";
				when "000011101001101100" => data <= "000000";
				when "000011101001101101" => data <= "000000";
				when "000011101001101110" => data <= "000000";
				when "000011101001101111" => data <= "000000";
				when "000011101001110000" => data <= "000000";
				when "000011101001110001" => data <= "000000";
				when "000011101001110010" => data <= "000000";
				when "000011101001110011" => data <= "000000";
				when "000011101001110100" => data <= "000000";
				when "000011101001110101" => data <= "000000";
				when "000011101001110110" => data <= "000000";
				when "000011101001110111" => data <= "000000";
				when "000011101001111000" => data <= "000000";
				when "000011101001111001" => data <= "000000";
				when "000011101001111010" => data <= "000000";
				when "000011101001111011" => data <= "000000";
				when "000011101001111100" => data <= "000000";
				when "000011101001111101" => data <= "000000";
				when "000011101001111110" => data <= "000000";
				when "000011101001111111" => data <= "000000";
				when "000011101010000000" => data <= "000000";
				when "000011101010000001" => data <= "000000";
				when "000011101010000010" => data <= "000000";
				when "000011101010000011" => data <= "000000";
				when "000011101010000100" => data <= "000000";
				when "000011101010000101" => data <= "000000";
				when "000011101010000110" => data <= "000000";
				when "000011101010000111" => data <= "000000";
				when "000011101010001000" => data <= "000000";
				when "000011101010001001" => data <= "000000";
				when "000011101010001010" => data <= "000000";
				when "000011101010001011" => data <= "000000";
				when "000011101010001100" => data <= "000000";
				when "000011101010001101" => data <= "000000";
				when "000011101010001110" => data <= "000000";
				when "000011101010001111" => data <= "000000";
				when "000011101010010000" => data <= "000000";
				when "000011101010010001" => data <= "000000";
				when "000011101010010010" => data <= "000000";
				when "000011101010010011" => data <= "000000";
				when "000011101010010100" => data <= "000000";
				when "000011101010010101" => data <= "000000";
				when "000011101010010110" => data <= "000000";
				when "000011101010010111" => data <= "000000";
				when "000011101010011000" => data <= "000000";
				when "000011101010011001" => data <= "000000";
				when "000011101010011010" => data <= "000000";
				when "000011101010011011" => data <= "000000";
				when "000011101010011100" => data <= "000000";
				when "000011101010011101" => data <= "000000";
				when "000011101010011110" => data <= "000000";
				when "000011101010011111" => data <= "000000";
				when "000011110000000000" => data <= "000000";
				when "000011110000000001" => data <= "000000";
				when "000011110000000010" => data <= "000000";
				when "000011110000000011" => data <= "000000";
				when "000011110000000100" => data <= "000000";
				when "000011110000000101" => data <= "000000";
				when "000011110000000110" => data <= "000000";
				when "000011110000000111" => data <= "000000";
				when "000011110000001000" => data <= "000000";
				when "000011110000001001" => data <= "000000";
				when "000011110000001010" => data <= "000000";
				when "000011110000001011" => data <= "000000";
				when "000011110000001100" => data <= "000000";
				when "000011110000001101" => data <= "000000";
				when "000011110000001110" => data <= "000000";
				when "000011110000001111" => data <= "000000";
				when "000011110000010000" => data <= "000000";
				when "000011110000010001" => data <= "000000";
				when "000011110000010010" => data <= "000000";
				when "000011110000010011" => data <= "000000";
				when "000011110000010100" => data <= "000000";
				when "000011110000010101" => data <= "000000";
				when "000011110000010110" => data <= "000000";
				when "000011110000010111" => data <= "000000";
				when "000011110000011000" => data <= "000000";
				when "000011110000011001" => data <= "000000";
				when "000011110000011010" => data <= "000000";
				when "000011110000011011" => data <= "000000";
				when "000011110000011100" => data <= "000000";
				when "000011110000011101" => data <= "000000";
				when "000011110000011110" => data <= "000000";
				when "000011110000011111" => data <= "000000";
				when "000011110000100000" => data <= "000000";
				when "000011110000100001" => data <= "000000";
				when "000011110000100010" => data <= "000000";
				when "000011110000100011" => data <= "000000";
				when "000011110000100100" => data <= "000000";
				when "000011110000100101" => data <= "000000";
				when "000011110000100110" => data <= "000000";
				when "000011110000100111" => data <= "000000";
				when "000011110000101000" => data <= "000000";
				when "000011110000101001" => data <= "000000";
				when "000011110000101010" => data <= "000000";
				when "000011110000101011" => data <= "000000";
				when "000011110000101100" => data <= "000000";
				when "000011110000101101" => data <= "000000";
				when "000011110000101110" => data <= "000000";
				when "000011110000101111" => data <= "000000";
				when "000011110000110000" => data <= "000000";
				when "000011110000110001" => data <= "000000";
				when "000011110000110010" => data <= "000000";
				when "000011110000110011" => data <= "000000";
				when "000011110000110100" => data <= "000000";
				when "000011110000110101" => data <= "000000";
				when "000011110000110110" => data <= "000000";
				when "000011110000110111" => data <= "000000";
				when "000011110000111000" => data <= "000000";
				when "000011110000111001" => data <= "000000";
				when "000011110000111010" => data <= "000000";
				when "000011110000111011" => data <= "000000";
				when "000011110000111100" => data <= "000000";
				when "000011110000111101" => data <= "000000";
				when "000011110000111110" => data <= "000000";
				when "000011110000111111" => data <= "000000";
				when "000011110001000000" => data <= "000000";
				when "000011110001000001" => data <= "000000";
				when "000011110001000010" => data <= "000000";
				when "000011110001000011" => data <= "000000";
				when "000011110001000100" => data <= "000000";
				when "000011110001000101" => data <= "000000";
				when "000011110001000110" => data <= "000000";
				when "000011110001000111" => data <= "000000";
				when "000011110001001000" => data <= "000000";
				when "000011110001001001" => data <= "000000";
				when "000011110001001010" => data <= "000000";
				when "000011110001001011" => data <= "000000";
				when "000011110001001100" => data <= "000000";
				when "000011110001001101" => data <= "000000";
				when "000011110001001110" => data <= "000000";
				when "000011110001001111" => data <= "000000";
				when "000011110001010000" => data <= "000000";
				when "000011110001010001" => data <= "000000";
				when "000011110001010010" => data <= "000000";
				when "000011110001010011" => data <= "000000";
				when "000011110001010100" => data <= "000000";
				when "000011110001010101" => data <= "000000";
				when "000011110001010110" => data <= "000000";
				when "000011110001010111" => data <= "000000";
				when "000011110001011000" => data <= "000000";
				when "000011110001011001" => data <= "000000";
				when "000011110001011010" => data <= "000000";
				when "000011110001011011" => data <= "000000";
				when "000011110001011100" => data <= "000000";
				when "000011110001011101" => data <= "000000";
				when "000011110001011110" => data <= "000000";
				when "000011110001011111" => data <= "000000";
				when "000011110001100000" => data <= "000000";
				when "000011110001100001" => data <= "000000";
				when "000011110001100010" => data <= "000000";
				when "000011110001100011" => data <= "000000";
				when "000011110001100100" => data <= "000000";
				when "000011110001100101" => data <= "000000";
				when "000011110001100110" => data <= "000000";
				when "000011110001100111" => data <= "000000";
				when "000011110001101000" => data <= "000000";
				when "000011110001101001" => data <= "000000";
				when "000011110001101010" => data <= "000000";
				when "000011110001101011" => data <= "000000";
				when "000011110001101100" => data <= "000000";
				when "000011110001101101" => data <= "000000";
				when "000011110001101110" => data <= "000000";
				when "000011110001101111" => data <= "000000";
				when "000011110001110000" => data <= "000000";
				when "000011110001110001" => data <= "000000";
				when "000011110001110010" => data <= "000000";
				when "000011110001110011" => data <= "000000";
				when "000011110001110100" => data <= "000000";
				when "000011110001110101" => data <= "000000";
				when "000011110001110110" => data <= "000000";
				when "000011110001110111" => data <= "000000";
				when "000011110001111000" => data <= "000000";
				when "000011110001111001" => data <= "000000";
				when "000011110001111010" => data <= "000000";
				when "000011110001111011" => data <= "000000";
				when "000011110001111100" => data <= "000000";
				when "000011110001111101" => data <= "000000";
				when "000011110001111110" => data <= "000000";
				when "000011110001111111" => data <= "000000";
				when "000011110010000000" => data <= "000000";
				when "000011110010000001" => data <= "000000";
				when "000011110010000010" => data <= "000000";
				when "000011110010000011" => data <= "000000";
				when "000011110010000100" => data <= "000000";
				when "000011110010000101" => data <= "000000";
				when "000011110010000110" => data <= "000000";
				when "000011110010000111" => data <= "000000";
				when "000011110010001000" => data <= "000000";
				when "000011110010001001" => data <= "000000";
				when "000011110010001010" => data <= "000000";
				when "000011110010001011" => data <= "000000";
				when "000011110010001100" => data <= "000000";
				when "000011110010001101" => data <= "000000";
				when "000011110010001110" => data <= "000000";
				when "000011110010001111" => data <= "000000";
				when "000011110010010000" => data <= "000000";
				when "000011110010010001" => data <= "000000";
				when "000011110010010010" => data <= "000000";
				when "000011110010010011" => data <= "000000";
				when "000011110010010100" => data <= "000000";
				when "000011110010010101" => data <= "000000";
				when "000011110010010110" => data <= "000000";
				when "000011110010010111" => data <= "000000";
				when "000011110010011000" => data <= "000000";
				when "000011110010011001" => data <= "000000";
				when "000011110010011010" => data <= "000000";
				when "000011110010011011" => data <= "000000";
				when "000011110010011100" => data <= "000000";
				when "000011110010011101" => data <= "000000";
				when "000011110010011110" => data <= "000000";
				when "000011110010011111" => data <= "000000";
				when "000011111000000000" => data <= "000000";
				when "000011111000000001" => data <= "000000";
				when "000011111000000010" => data <= "000000";
				when "000011111000000011" => data <= "000000";
				when "000011111000000100" => data <= "000000";
				when "000011111000000101" => data <= "000000";
				when "000011111000000110" => data <= "000000";
				when "000011111000000111" => data <= "000000";
				when "000011111000001000" => data <= "000000";
				when "000011111000001001" => data <= "000000";
				when "000011111000001010" => data <= "000000";
				when "000011111000001011" => data <= "000000";
				when "000011111000001100" => data <= "000000";
				when "000011111000001101" => data <= "000000";
				when "000011111000001110" => data <= "000000";
				when "000011111000001111" => data <= "000000";
				when "000011111000010000" => data <= "000000";
				when "000011111000010001" => data <= "000000";
				when "000011111000010010" => data <= "000000";
				when "000011111000010011" => data <= "000000";
				when "000011111000010100" => data <= "000000";
				when "000011111000010101" => data <= "000000";
				when "000011111000010110" => data <= "000000";
				when "000011111000010111" => data <= "000000";
				when "000011111000011000" => data <= "000000";
				when "000011111000011001" => data <= "000000";
				when "000011111000011010" => data <= "000000";
				when "000011111000011011" => data <= "000000";
				when "000011111000011100" => data <= "000000";
				when "000011111000011101" => data <= "000000";
				when "000011111000011110" => data <= "000000";
				when "000011111000011111" => data <= "000000";
				when "000011111000100000" => data <= "000000";
				when "000011111000100001" => data <= "000000";
				when "000011111000100010" => data <= "000000";
				when "000011111000100011" => data <= "000000";
				when "000011111000100100" => data <= "000000";
				when "000011111000100101" => data <= "000000";
				when "000011111000100110" => data <= "000000";
				when "000011111000100111" => data <= "000000";
				when "000011111000101000" => data <= "000000";
				when "000011111000101001" => data <= "000000";
				when "000011111000101010" => data <= "000000";
				when "000011111000101011" => data <= "000000";
				when "000011111000101100" => data <= "000000";
				when "000011111000101101" => data <= "000000";
				when "000011111000101110" => data <= "000000";
				when "000011111000101111" => data <= "000000";
				when "000011111000110000" => data <= "000000";
				when "000011111000110001" => data <= "000000";
				when "000011111000110010" => data <= "000000";
				when "000011111000110011" => data <= "000000";
				when "000011111000110100" => data <= "000000";
				when "000011111000110101" => data <= "000000";
				when "000011111000110110" => data <= "000000";
				when "000011111000110111" => data <= "000000";
				when "000011111000111000" => data <= "000000";
				when "000011111000111001" => data <= "000000";
				when "000011111000111010" => data <= "000000";
				when "000011111000111011" => data <= "000000";
				when "000011111000111100" => data <= "000000";
				when "000011111000111101" => data <= "000000";
				when "000011111000111110" => data <= "000000";
				when "000011111000111111" => data <= "000000";
				when "000011111001000000" => data <= "000000";
				when "000011111001000001" => data <= "000000";
				when "000011111001000010" => data <= "000000";
				when "000011111001000011" => data <= "000000";
				when "000011111001000100" => data <= "000000";
				when "000011111001000101" => data <= "000000";
				when "000011111001000110" => data <= "000000";
				when "000011111001000111" => data <= "000000";
				when "000011111001001000" => data <= "000000";
				when "000011111001001001" => data <= "000000";
				when "000011111001001010" => data <= "000000";
				when "000011111001001011" => data <= "000000";
				when "000011111001001100" => data <= "000000";
				when "000011111001001101" => data <= "000000";
				when "000011111001001110" => data <= "000000";
				when "000011111001001111" => data <= "000000";
				when "000011111001010000" => data <= "000000";
				when "000011111001010001" => data <= "000000";
				when "000011111001010010" => data <= "000000";
				when "000011111001010011" => data <= "000000";
				when "000011111001010100" => data <= "000000";
				when "000011111001010101" => data <= "000000";
				when "000011111001010110" => data <= "000000";
				when "000011111001010111" => data <= "000000";
				when "000011111001011000" => data <= "000000";
				when "000011111001011001" => data <= "000000";
				when "000011111001011010" => data <= "000000";
				when "000011111001011011" => data <= "000000";
				when "000011111001011100" => data <= "000000";
				when "000011111001011101" => data <= "000000";
				when "000011111001011110" => data <= "000000";
				when "000011111001011111" => data <= "000000";
				when "000011111001100000" => data <= "000000";
				when "000011111001100001" => data <= "000000";
				when "000011111001100010" => data <= "000000";
				when "000011111001100011" => data <= "000000";
				when "000011111001100100" => data <= "000000";
				when "000011111001100101" => data <= "000000";
				when "000011111001100110" => data <= "000000";
				when "000011111001100111" => data <= "000000";
				when "000011111001101000" => data <= "000000";
				when "000011111001101001" => data <= "000000";
				when "000011111001101010" => data <= "000000";
				when "000011111001101011" => data <= "000000";
				when "000011111001101100" => data <= "000000";
				when "000011111001101101" => data <= "000000";
				when "000011111001101110" => data <= "000000";
				when "000011111001101111" => data <= "000000";
				when "000011111001110000" => data <= "000000";
				when "000011111001110001" => data <= "000000";
				when "000011111001110010" => data <= "000000";
				when "000011111001110011" => data <= "000000";
				when "000011111001110100" => data <= "000000";
				when "000011111001110101" => data <= "000000";
				when "000011111001110110" => data <= "000000";
				when "000011111001110111" => data <= "000000";
				when "000011111001111000" => data <= "000000";
				when "000011111001111001" => data <= "000000";
				when "000011111001111010" => data <= "000000";
				when "000011111001111011" => data <= "000000";
				when "000011111001111100" => data <= "000000";
				when "000011111001111101" => data <= "000000";
				when "000011111001111110" => data <= "000000";
				when "000011111001111111" => data <= "000000";
				when "000011111010000000" => data <= "000000";
				when "000011111010000001" => data <= "000000";
				when "000011111010000010" => data <= "000000";
				when "000011111010000011" => data <= "000000";
				when "000011111010000100" => data <= "000000";
				when "000011111010000101" => data <= "000000";
				when "000011111010000110" => data <= "000000";
				when "000011111010000111" => data <= "000000";
				when "000011111010001000" => data <= "000000";
				when "000011111010001001" => data <= "000000";
				when "000011111010001010" => data <= "000000";
				when "000011111010001011" => data <= "000000";
				when "000011111010001100" => data <= "000000";
				when "000011111010001101" => data <= "000000";
				when "000011111010001110" => data <= "000000";
				when "000011111010001111" => data <= "000000";
				when "000011111010010000" => data <= "000000";
				when "000011111010010001" => data <= "000000";
				when "000011111010010010" => data <= "000000";
				when "000011111010010011" => data <= "000000";
				when "000011111010010100" => data <= "000000";
				when "000011111010010101" => data <= "000000";
				when "000011111010010110" => data <= "000000";
				when "000011111010010111" => data <= "000000";
				when "000011111010011000" => data <= "000000";
				when "000011111010011001" => data <= "000000";
				when "000011111010011010" => data <= "000000";
				when "000011111010011011" => data <= "000000";
				when "000011111010011100" => data <= "000000";
				when "000011111010011101" => data <= "000000";
				when "000011111010011110" => data <= "000000";
				when "000011111010011111" => data <= "000000";
				when "000100000000000000" => data <= "000000";
				when "000100000000000001" => data <= "000000";
				when "000100000000000010" => data <= "000000";
				when "000100000000000011" => data <= "000000";
				when "000100000000000100" => data <= "000000";
				when "000100000000000101" => data <= "000000";
				when "000100000000000110" => data <= "000000";
				when "000100000000000111" => data <= "000000";
				when "000100000000001000" => data <= "000000";
				when "000100000000001001" => data <= "000000";
				when "000100000000001010" => data <= "000000";
				when "000100000000001011" => data <= "000000";
				when "000100000000001100" => data <= "000000";
				when "000100000000001101" => data <= "000000";
				when "000100000000001110" => data <= "000000";
				when "000100000000001111" => data <= "000000";
				when "000100000000010000" => data <= "000000";
				when "000100000000010001" => data <= "000000";
				when "000100000000010010" => data <= "000000";
				when "000100000000010011" => data <= "000000";
				when "000100000000010100" => data <= "000000";
				when "000100000000010101" => data <= "000000";
				when "000100000000010110" => data <= "000000";
				when "000100000000010111" => data <= "000000";
				when "000100000000011000" => data <= "000000";
				when "000100000000011001" => data <= "000000";
				when "000100000000011010" => data <= "000000";
				when "000100000000011011" => data <= "000000";
				when "000100000000011100" => data <= "000000";
				when "000100000000011101" => data <= "000000";
				when "000100000000011110" => data <= "000000";
				when "000100000000011111" => data <= "000000";
				when "000100000000100000" => data <= "000000";
				when "000100000000100001" => data <= "000000";
				when "000100000000100010" => data <= "000000";
				when "000100000000100011" => data <= "000000";
				when "000100000000100100" => data <= "000000";
				when "000100000000100101" => data <= "000000";
				when "000100000000100110" => data <= "000000";
				when "000100000000100111" => data <= "000000";
				when "000100000000101000" => data <= "000000";
				when "000100000000101001" => data <= "000000";
				when "000100000000101010" => data <= "000000";
				when "000100000000101011" => data <= "000000";
				when "000100000000101100" => data <= "000000";
				when "000100000000101101" => data <= "000000";
				when "000100000000101110" => data <= "000000";
				when "000100000000101111" => data <= "000000";
				when "000100000000110000" => data <= "000000";
				when "000100000000110001" => data <= "000000";
				when "000100000000110010" => data <= "000000";
				when "000100000000110011" => data <= "000000";
				when "000100000000110100" => data <= "000000";
				when "000100000000110101" => data <= "000000";
				when "000100000000110110" => data <= "000000";
				when "000100000000110111" => data <= "000000";
				when "000100000000111000" => data <= "000000";
				when "000100000000111001" => data <= "000000";
				when "000100000000111010" => data <= "000000";
				when "000100000000111011" => data <= "000000";
				when "000100000000111100" => data <= "000000";
				when "000100000000111101" => data <= "000000";
				when "000100000000111110" => data <= "000000";
				when "000100000000111111" => data <= "000000";
				when "000100000001000000" => data <= "000000";
				when "000100000001000001" => data <= "000000";
				when "000100000001000010" => data <= "000000";
				when "000100000001000011" => data <= "000000";
				when "000100000001000100" => data <= "000000";
				when "000100000001000101" => data <= "000000";
				when "000100000001000110" => data <= "000000";
				when "000100000001000111" => data <= "000000";
				when "000100000001001000" => data <= "000000";
				when "000100000001001001" => data <= "000000";
				when "000100000001001010" => data <= "000000";
				when "000100000001001011" => data <= "000000";
				when "000100000001001100" => data <= "000000";
				when "000100000001001101" => data <= "000000";
				when "000100000001001110" => data <= "000000";
				when "000100000001001111" => data <= "000000";
				when "000100000001010000" => data <= "000000";
				when "000100000001010001" => data <= "000000";
				when "000100000001010010" => data <= "000000";
				when "000100000001010011" => data <= "000000";
				when "000100000001010100" => data <= "000000";
				when "000100000001010101" => data <= "000000";
				when "000100000001010110" => data <= "000000";
				when "000100000001010111" => data <= "000000";
				when "000100000001011000" => data <= "000000";
				when "000100000001011001" => data <= "000000";
				when "000100000001011010" => data <= "000000";
				when "000100000001011011" => data <= "000000";
				when "000100000001011100" => data <= "000000";
				when "000100000001011101" => data <= "000000";
				when "000100000001011110" => data <= "000000";
				when "000100000001011111" => data <= "000000";
				when "000100000001100000" => data <= "000000";
				when "000100000001100001" => data <= "000000";
				when "000100000001100010" => data <= "000000";
				when "000100000001100011" => data <= "000000";
				when "000100000001100100" => data <= "000000";
				when "000100000001100101" => data <= "000000";
				when "000100000001100110" => data <= "000000";
				when "000100000001100111" => data <= "000000";
				when "000100000001101000" => data <= "000000";
				when "000100000001101001" => data <= "000000";
				when "000100000001101010" => data <= "000000";
				when "000100000001101011" => data <= "000000";
				when "000100000001101100" => data <= "000000";
				when "000100000001101101" => data <= "000000";
				when "000100000001101110" => data <= "000000";
				when "000100000001101111" => data <= "000000";
				when "000100000001110000" => data <= "000000";
				when "000100000001110001" => data <= "000000";
				when "000100000001110010" => data <= "000000";
				when "000100000001110011" => data <= "000000";
				when "000100000001110100" => data <= "000000";
				when "000100000001110101" => data <= "000000";
				when "000100000001110110" => data <= "000000";
				when "000100000001110111" => data <= "000000";
				when "000100000001111000" => data <= "000000";
				when "000100000001111001" => data <= "000000";
				when "000100000001111010" => data <= "000000";
				when "000100000001111011" => data <= "000000";
				when "000100000001111100" => data <= "000000";
				when "000100000001111101" => data <= "000000";
				when "000100000001111110" => data <= "000000";
				when "000100000001111111" => data <= "000000";
				when "000100000010000000" => data <= "000000";
				when "000100000010000001" => data <= "000000";
				when "000100000010000010" => data <= "000000";
				when "000100000010000011" => data <= "000000";
				when "000100000010000100" => data <= "000000";
				when "000100000010000101" => data <= "000000";
				when "000100000010000110" => data <= "000000";
				when "000100000010000111" => data <= "000000";
				when "000100000010001000" => data <= "000000";
				when "000100000010001001" => data <= "000000";
				when "000100000010001010" => data <= "000000";
				when "000100000010001011" => data <= "000000";
				when "000100000010001100" => data <= "000000";
				when "000100000010001101" => data <= "000000";
				when "000100000010001110" => data <= "000000";
				when "000100000010001111" => data <= "000000";
				when "000100000010010000" => data <= "000000";
				when "000100000010010001" => data <= "000000";
				when "000100000010010010" => data <= "000000";
				when "000100000010010011" => data <= "000000";
				when "000100000010010100" => data <= "000000";
				when "000100000010010101" => data <= "000000";
				when "000100000010010110" => data <= "000000";
				when "000100000010010111" => data <= "000000";
				when "000100000010011000" => data <= "000000";
				when "000100000010011001" => data <= "000000";
				when "000100000010011010" => data <= "000000";
				when "000100000010011011" => data <= "000000";
				when "000100000010011100" => data <= "000000";
				when "000100000010011101" => data <= "000000";
				when "000100000010011110" => data <= "000000";
				when "000100000010011111" => data <= "000000";
				when "000100001000000000" => data <= "000000";
				when "000100001000000001" => data <= "000000";
				when "000100001000000010" => data <= "000000";
				when "000100001000000011" => data <= "000000";
				when "000100001000000100" => data <= "000000";
				when "000100001000000101" => data <= "000000";
				when "000100001000000110" => data <= "000000";
				when "000100001000000111" => data <= "000000";
				when "000100001000001000" => data <= "000000";
				when "000100001000001001" => data <= "000000";
				when "000100001000001010" => data <= "000000";
				when "000100001000001011" => data <= "000000";
				when "000100001000001100" => data <= "000000";
				when "000100001000001101" => data <= "000000";
				when "000100001000001110" => data <= "000000";
				when "000100001000001111" => data <= "000000";
				when "000100001000010000" => data <= "000000";
				when "000100001000010001" => data <= "000000";
				when "000100001000010010" => data <= "000000";
				when "000100001000010011" => data <= "000000";
				when "000100001000010100" => data <= "000000";
				when "000100001000010101" => data <= "000000";
				when "000100001000010110" => data <= "000000";
				when "000100001000010111" => data <= "000000";
				when "000100001000011000" => data <= "000000";
				when "000100001000011001" => data <= "000000";
				when "000100001000011010" => data <= "000000";
				when "000100001000011011" => data <= "000000";
				when "000100001000011100" => data <= "000000";
				when "000100001000011101" => data <= "000000";
				when "000100001000011110" => data <= "000000";
				when "000100001000011111" => data <= "000000";
				when "000100001000100000" => data <= "000000";
				when "000100001000100001" => data <= "000000";
				when "000100001000100010" => data <= "000000";
				when "000100001000100011" => data <= "000000";
				when "000100001000100100" => data <= "000000";
				when "000100001000100101" => data <= "000000";
				when "000100001000100110" => data <= "000000";
				when "000100001000100111" => data <= "000000";
				when "000100001000101000" => data <= "000000";
				when "000100001000101001" => data <= "000000";
				when "000100001000101010" => data <= "000000";
				when "000100001000101011" => data <= "000000";
				when "000100001000101100" => data <= "000000";
				when "000100001000101101" => data <= "000000";
				when "000100001000101110" => data <= "000000";
				when "000100001000101111" => data <= "000000";
				when "000100001000110000" => data <= "000000";
				when "000100001000110001" => data <= "000000";
				when "000100001000110010" => data <= "000000";
				when "000100001000110011" => data <= "000000";
				when "000100001000110100" => data <= "000000";
				when "000100001000110101" => data <= "000000";
				when "000100001000110110" => data <= "000000";
				when "000100001000110111" => data <= "000000";
				when "000100001000111000" => data <= "000000";
				when "000100001000111001" => data <= "000000";
				when "000100001000111010" => data <= "000000";
				when "000100001000111011" => data <= "000000";
				when "000100001000111100" => data <= "000000";
				when "000100001000111101" => data <= "000000";
				when "000100001000111110" => data <= "000000";
				when "000100001000111111" => data <= "000000";
				when "000100001001000000" => data <= "000000";
				when "000100001001000001" => data <= "000000";
				when "000100001001000010" => data <= "000000";
				when "000100001001000011" => data <= "000000";
				when "000100001001000100" => data <= "000000";
				when "000100001001000101" => data <= "000000";
				when "000100001001000110" => data <= "000000";
				when "000100001001000111" => data <= "000000";
				when "000100001001001000" => data <= "000000";
				when "000100001001001001" => data <= "000000";
				when "000100001001001010" => data <= "000000";
				when "000100001001001011" => data <= "000000";
				when "000100001001001100" => data <= "000000";
				when "000100001001001101" => data <= "000000";
				when "000100001001001110" => data <= "000000";
				when "000100001001001111" => data <= "000000";
				when "000100001001010000" => data <= "000000";
				when "000100001001010001" => data <= "000000";
				when "000100001001010010" => data <= "000000";
				when "000100001001010011" => data <= "000000";
				when "000100001001010100" => data <= "000000";
				when "000100001001010101" => data <= "000000";
				when "000100001001010110" => data <= "000000";
				when "000100001001010111" => data <= "000000";
				when "000100001001011000" => data <= "000000";
				when "000100001001011001" => data <= "000000";
				when "000100001001011010" => data <= "000000";
				when "000100001001011011" => data <= "000000";
				when "000100001001011100" => data <= "000000";
				when "000100001001011101" => data <= "000000";
				when "000100001001011110" => data <= "000000";
				when "000100001001011111" => data <= "000000";
				when "000100001001100000" => data <= "000000";
				when "000100001001100001" => data <= "000000";
				when "000100001001100010" => data <= "000000";
				when "000100001001100011" => data <= "000000";
				when "000100001001100100" => data <= "000000";
				when "000100001001100101" => data <= "000000";
				when "000100001001100110" => data <= "000000";
				when "000100001001100111" => data <= "000000";
				when "000100001001101000" => data <= "000000";
				when "000100001001101001" => data <= "000000";
				when "000100001001101010" => data <= "000000";
				when "000100001001101011" => data <= "000000";
				when "000100001001101100" => data <= "000000";
				when "000100001001101101" => data <= "000000";
				when "000100001001101110" => data <= "000000";
				when "000100001001101111" => data <= "000000";
				when "000100001001110000" => data <= "000000";
				when "000100001001110001" => data <= "000000";
				when "000100001001110010" => data <= "000000";
				when "000100001001110011" => data <= "000000";
				when "000100001001110100" => data <= "000000";
				when "000100001001110101" => data <= "000000";
				when "000100001001110110" => data <= "000000";
				when "000100001001110111" => data <= "000000";
				when "000100001001111000" => data <= "000000";
				when "000100001001111001" => data <= "000000";
				when "000100001001111010" => data <= "000000";
				when "000100001001111011" => data <= "000000";
				when "000100001001111100" => data <= "000000";
				when "000100001001111101" => data <= "000000";
				when "000100001001111110" => data <= "000000";
				when "000100001001111111" => data <= "000000";
				when "000100001010000000" => data <= "000000";
				when "000100001010000001" => data <= "000000";
				when "000100001010000010" => data <= "000000";
				when "000100001010000011" => data <= "000000";
				when "000100001010000100" => data <= "000000";
				when "000100001010000101" => data <= "000000";
				when "000100001010000110" => data <= "000000";
				when "000100001010000111" => data <= "000000";
				when "000100001010001000" => data <= "000000";
				when "000100001010001001" => data <= "000000";
				when "000100001010001010" => data <= "000000";
				when "000100001010001011" => data <= "000000";
				when "000100001010001100" => data <= "000000";
				when "000100001010001101" => data <= "000000";
				when "000100001010001110" => data <= "000000";
				when "000100001010001111" => data <= "000000";
				when "000100001010010000" => data <= "000000";
				when "000100001010010001" => data <= "000000";
				when "000100001010010010" => data <= "000000";
				when "000100001010010011" => data <= "000000";
				when "000100001010010100" => data <= "000000";
				when "000100001010010101" => data <= "000000";
				when "000100001010010110" => data <= "000000";
				when "000100001010010111" => data <= "000000";
				when "000100001010011000" => data <= "000000";
				when "000100001010011001" => data <= "000000";
				when "000100001010011010" => data <= "000000";
				when "000100001010011011" => data <= "000000";
				when "000100001010011100" => data <= "000000";
				when "000100001010011101" => data <= "000000";
				when "000100001010011110" => data <= "000000";
				when "000100001010011111" => data <= "000000";
				when "000100010000000000" => data <= "000000";
				when "000100010000000001" => data <= "000000";
				when "000100010000000010" => data <= "000000";
				when "000100010000000011" => data <= "000000";
				when "000100010000000100" => data <= "000000";
				when "000100010000000101" => data <= "000000";
				when "000100010000000110" => data <= "000000";
				when "000100010000000111" => data <= "000000";
				when "000100010000001000" => data <= "000000";
				when "000100010000001001" => data <= "000000";
				when "000100010000001010" => data <= "000000";
				when "000100010000001011" => data <= "000000";
				when "000100010000001100" => data <= "000000";
				when "000100010000001101" => data <= "000000";
				when "000100010000001110" => data <= "000000";
				when "000100010000001111" => data <= "000000";
				when "000100010000010000" => data <= "000000";
				when "000100010000010001" => data <= "000000";
				when "000100010000010010" => data <= "000000";
				when "000100010000010011" => data <= "000000";
				when "000100010000010100" => data <= "000000";
				when "000100010000010101" => data <= "000000";
				when "000100010000010110" => data <= "000000";
				when "000100010000010111" => data <= "000000";
				when "000100010000011000" => data <= "000000";
				when "000100010000011001" => data <= "000000";
				when "000100010000011010" => data <= "000000";
				when "000100010000011011" => data <= "000000";
				when "000100010000011100" => data <= "000000";
				when "000100010000011101" => data <= "000000";
				when "000100010000011110" => data <= "000000";
				when "000100010000011111" => data <= "000000";
				when "000100010000100000" => data <= "000000";
				when "000100010000100001" => data <= "000000";
				when "000100010000100010" => data <= "000000";
				when "000100010000100011" => data <= "000000";
				when "000100010000100100" => data <= "000000";
				when "000100010000100101" => data <= "000000";
				when "000100010000100110" => data <= "000000";
				when "000100010000100111" => data <= "000000";
				when "000100010000101000" => data <= "000000";
				when "000100010000101001" => data <= "000000";
				when "000100010000101010" => data <= "000000";
				when "000100010000101011" => data <= "000000";
				when "000100010000101100" => data <= "000000";
				when "000100010000101101" => data <= "000000";
				when "000100010000101110" => data <= "000000";
				when "000100010000101111" => data <= "000000";
				when "000100010000110000" => data <= "000000";
				when "000100010000110001" => data <= "000000";
				when "000100010000110010" => data <= "000000";
				when "000100010000110011" => data <= "000000";
				when "000100010000110100" => data <= "000000";
				when "000100010000110101" => data <= "000000";
				when "000100010000110110" => data <= "000000";
				when "000100010000110111" => data <= "000000";
				when "000100010000111000" => data <= "000000";
				when "000100010000111001" => data <= "000000";
				when "000100010000111010" => data <= "000000";
				when "000100010000111011" => data <= "000000";
				when "000100010000111100" => data <= "000000";
				when "000100010000111101" => data <= "000000";
				when "000100010000111110" => data <= "000000";
				when "000100010000111111" => data <= "000000";
				when "000100010001000000" => data <= "000000";
				when "000100010001000001" => data <= "000000";
				when "000100010001000010" => data <= "000000";
				when "000100010001000011" => data <= "000000";
				when "000100010001000100" => data <= "000000";
				when "000100010001000101" => data <= "000000";
				when "000100010001000110" => data <= "000000";
				when "000100010001000111" => data <= "000000";
				when "000100010001001000" => data <= "000000";
				when "000100010001001001" => data <= "000000";
				when "000100010001001010" => data <= "000000";
				when "000100010001001011" => data <= "000000";
				when "000100010001001100" => data <= "000000";
				when "000100010001001101" => data <= "000000";
				when "000100010001001110" => data <= "000000";
				when "000100010001001111" => data <= "000000";
				when "000100010001010000" => data <= "000000";
				when "000100010001010001" => data <= "000000";
				when "000100010001010010" => data <= "000000";
				when "000100010001010011" => data <= "000000";
				when "000100010001010100" => data <= "000000";
				when "000100010001010101" => data <= "000000";
				when "000100010001010110" => data <= "000000";
				when "000100010001010111" => data <= "000000";
				when "000100010001011000" => data <= "000000";
				when "000100010001011001" => data <= "000000";
				when "000100010001011010" => data <= "000000";
				when "000100010001011011" => data <= "000000";
				when "000100010001011100" => data <= "000000";
				when "000100010001011101" => data <= "000000";
				when "000100010001011110" => data <= "000000";
				when "000100010001011111" => data <= "000000";
				when "000100010001100000" => data <= "000000";
				when "000100010001100001" => data <= "000000";
				when "000100010001100010" => data <= "000000";
				when "000100010001100011" => data <= "000000";
				when "000100010001100100" => data <= "000000";
				when "000100010001100101" => data <= "000000";
				when "000100010001100110" => data <= "000000";
				when "000100010001100111" => data <= "000000";
				when "000100010001101000" => data <= "000000";
				when "000100010001101001" => data <= "000000";
				when "000100010001101010" => data <= "000000";
				when "000100010001101011" => data <= "000000";
				when "000100010001101100" => data <= "000000";
				when "000100010001101101" => data <= "000000";
				when "000100010001101110" => data <= "000000";
				when "000100010001101111" => data <= "000000";
				when "000100010001110000" => data <= "000000";
				when "000100010001110001" => data <= "000000";
				when "000100010001110010" => data <= "000000";
				when "000100010001110011" => data <= "000000";
				when "000100010001110100" => data <= "000000";
				when "000100010001110101" => data <= "000000";
				when "000100010001110110" => data <= "000000";
				when "000100010001110111" => data <= "000000";
				when "000100010001111000" => data <= "000000";
				when "000100010001111001" => data <= "000000";
				when "000100010001111010" => data <= "000000";
				when "000100010001111011" => data <= "000000";
				when "000100010001111100" => data <= "000000";
				when "000100010001111101" => data <= "000000";
				when "000100010001111110" => data <= "000000";
				when "000100010001111111" => data <= "000000";
				when "000100010010000000" => data <= "000000";
				when "000100010010000001" => data <= "000000";
				when "000100010010000010" => data <= "000000";
				when "000100010010000011" => data <= "000000";
				when "000100010010000100" => data <= "000000";
				when "000100010010000101" => data <= "000000";
				when "000100010010000110" => data <= "000000";
				when "000100010010000111" => data <= "000000";
				when "000100010010001000" => data <= "000000";
				when "000100010010001001" => data <= "000000";
				when "000100010010001010" => data <= "000000";
				when "000100010010001011" => data <= "000000";
				when "000100010010001100" => data <= "000000";
				when "000100010010001101" => data <= "000000";
				when "000100010010001110" => data <= "000000";
				when "000100010010001111" => data <= "000000";
				when "000100010010010000" => data <= "000000";
				when "000100010010010001" => data <= "000000";
				when "000100010010010010" => data <= "000000";
				when "000100010010010011" => data <= "000000";
				when "000100010010010100" => data <= "000000";
				when "000100010010010101" => data <= "000000";
				when "000100010010010110" => data <= "000000";
				when "000100010010010111" => data <= "000000";
				when "000100010010011000" => data <= "000000";
				when "000100010010011001" => data <= "000000";
				when "000100010010011010" => data <= "000000";
				when "000100010010011011" => data <= "000000";
				when "000100010010011100" => data <= "000000";
				when "000100010010011101" => data <= "000000";
				when "000100010010011110" => data <= "000000";
				when "000100010010011111" => data <= "000000";
				when "000100011000000000" => data <= "000000";
				when "000100011000000001" => data <= "000000";
				when "000100011000000010" => data <= "000000";
				when "000100011000000011" => data <= "000000";
				when "000100011000000100" => data <= "000000";
				when "000100011000000101" => data <= "000000";
				when "000100011000000110" => data <= "000000";
				when "000100011000000111" => data <= "000000";
				when "000100011000001000" => data <= "000000";
				when "000100011000001001" => data <= "000000";
				when "000100011000001010" => data <= "000000";
				when "000100011000001011" => data <= "000000";
				when "000100011000001100" => data <= "000000";
				when "000100011000001101" => data <= "000000";
				when "000100011000001110" => data <= "000000";
				when "000100011000001111" => data <= "000000";
				when "000100011000010000" => data <= "000000";
				when "000100011000010001" => data <= "000000";
				when "000100011000010010" => data <= "000000";
				when "000100011000010011" => data <= "000000";
				when "000100011000010100" => data <= "000000";
				when "000100011000010101" => data <= "000000";
				when "000100011000010110" => data <= "000000";
				when "000100011000010111" => data <= "000000";
				when "000100011000011000" => data <= "000000";
				when "000100011000011001" => data <= "000000";
				when "000100011000011010" => data <= "000000";
				when "000100011000011011" => data <= "000000";
				when "000100011000011100" => data <= "000000";
				when "000100011000011101" => data <= "000000";
				when "000100011000011110" => data <= "000000";
				when "000100011000011111" => data <= "000000";
				when "000100011000100000" => data <= "000000";
				when "000100011000100001" => data <= "000000";
				when "000100011000100010" => data <= "000000";
				when "000100011000100011" => data <= "000000";
				when "000100011000100100" => data <= "000000";
				when "000100011000100101" => data <= "000000";
				when "000100011000100110" => data <= "000000";
				when "000100011000100111" => data <= "000000";
				when "000100011000101000" => data <= "000000";
				when "000100011000101001" => data <= "000000";
				when "000100011000101010" => data <= "000000";
				when "000100011000101011" => data <= "000000";
				when "000100011000101100" => data <= "000000";
				when "000100011000101101" => data <= "000000";
				when "000100011000101110" => data <= "000000";
				when "000100011000101111" => data <= "000000";
				when "000100011000110000" => data <= "000000";
				when "000100011000110001" => data <= "000000";
				when "000100011000110010" => data <= "000000";
				when "000100011000110011" => data <= "000000";
				when "000100011000110100" => data <= "000000";
				when "000100011000110101" => data <= "000000";
				when "000100011000110110" => data <= "000000";
				when "000100011000110111" => data <= "000000";
				when "000100011000111000" => data <= "000000";
				when "000100011000111001" => data <= "000000";
				when "000100011000111010" => data <= "000000";
				when "000100011000111011" => data <= "000000";
				when "000100011000111100" => data <= "000000";
				when "000100011000111101" => data <= "000000";
				when "000100011000111110" => data <= "000000";
				when "000100011000111111" => data <= "000000";
				when "000100011001000000" => data <= "000000";
				when "000100011001000001" => data <= "000000";
				when "000100011001000010" => data <= "000000";
				when "000100011001000011" => data <= "000000";
				when "000100011001000100" => data <= "000000";
				when "000100011001000101" => data <= "000000";
				when "000100011001000110" => data <= "000000";
				when "000100011001000111" => data <= "000000";
				when "000100011001001000" => data <= "000000";
				when "000100011001001001" => data <= "000000";
				when "000100011001001010" => data <= "000000";
				when "000100011001001011" => data <= "000000";
				when "000100011001001100" => data <= "000000";
				when "000100011001001101" => data <= "000000";
				when "000100011001001110" => data <= "000000";
				when "000100011001001111" => data <= "000000";
				when "000100011001010000" => data <= "000000";
				when "000100011001010001" => data <= "000000";
				when "000100011001010010" => data <= "000000";
				when "000100011001010011" => data <= "000000";
				when "000100011001010100" => data <= "000000";
				when "000100011001010101" => data <= "000000";
				when "000100011001010110" => data <= "000000";
				when "000100011001010111" => data <= "000000";
				when "000100011001011000" => data <= "000000";
				when "000100011001011001" => data <= "000000";
				when "000100011001011010" => data <= "000000";
				when "000100011001011011" => data <= "000000";
				when "000100011001011100" => data <= "000000";
				when "000100011001011101" => data <= "000000";
				when "000100011001011110" => data <= "000000";
				when "000100011001011111" => data <= "000000";
				when "000100011001100000" => data <= "000000";
				when "000100011001100001" => data <= "000000";
				when "000100011001100010" => data <= "000000";
				when "000100011001100011" => data <= "000000";
				when "000100011001100100" => data <= "000000";
				when "000100011001100101" => data <= "000000";
				when "000100011001100110" => data <= "000000";
				when "000100011001100111" => data <= "000000";
				when "000100011001101000" => data <= "000000";
				when "000100011001101001" => data <= "000000";
				when "000100011001101010" => data <= "000000";
				when "000100011001101011" => data <= "000000";
				when "000100011001101100" => data <= "000000";
				when "000100011001101101" => data <= "000000";
				when "000100011001101110" => data <= "000000";
				when "000100011001101111" => data <= "000000";
				when "000100011001110000" => data <= "000000";
				when "000100011001110001" => data <= "000000";
				when "000100011001110010" => data <= "000000";
				when "000100011001110011" => data <= "000000";
				when "000100011001110100" => data <= "000000";
				when "000100011001110101" => data <= "000000";
				when "000100011001110110" => data <= "000000";
				when "000100011001110111" => data <= "000000";
				when "000100011001111000" => data <= "000000";
				when "000100011001111001" => data <= "000000";
				when "000100011001111010" => data <= "000000";
				when "000100011001111011" => data <= "000000";
				when "000100011001111100" => data <= "000000";
				when "000100011001111101" => data <= "000000";
				when "000100011001111110" => data <= "000000";
				when "000100011001111111" => data <= "000000";
				when "000100011010000000" => data <= "000000";
				when "000100011010000001" => data <= "000000";
				when "000100011010000010" => data <= "000000";
				when "000100011010000011" => data <= "000000";
				when "000100011010000100" => data <= "000000";
				when "000100011010000101" => data <= "000000";
				when "000100011010000110" => data <= "000000";
				when "000100011010000111" => data <= "000000";
				when "000100011010001000" => data <= "000000";
				when "000100011010001001" => data <= "000000";
				when "000100011010001010" => data <= "000000";
				when "000100011010001011" => data <= "000000";
				when "000100011010001100" => data <= "000000";
				when "000100011010001101" => data <= "000000";
				when "000100011010001110" => data <= "000000";
				when "000100011010001111" => data <= "000000";
				when "000100011010010000" => data <= "000000";
				when "000100011010010001" => data <= "000000";
				when "000100011010010010" => data <= "000000";
				when "000100011010010011" => data <= "000000";
				when "000100011010010100" => data <= "000000";
				when "000100011010010101" => data <= "000000";
				when "000100011010010110" => data <= "000000";
				when "000100011010010111" => data <= "000000";
				when "000100011010011000" => data <= "000000";
				when "000100011010011001" => data <= "000000";
				when "000100011010011010" => data <= "000000";
				when "000100011010011011" => data <= "000000";
				when "000100011010011100" => data <= "000000";
				when "000100011010011101" => data <= "000000";
				when "000100011010011110" => data <= "000000";
				when "000100011010011111" => data <= "000000";
				when "000100100000000000" => data <= "000000";
				when "000100100000000001" => data <= "000000";
				when "000100100000000010" => data <= "000000";
				when "000100100000000011" => data <= "000000";
				when "000100100000000100" => data <= "000000";
				when "000100100000000101" => data <= "000000";
				when "000100100000000110" => data <= "000000";
				when "000100100000000111" => data <= "000000";
				when "000100100000001000" => data <= "000000";
				when "000100100000001001" => data <= "000000";
				when "000100100000001010" => data <= "000000";
				when "000100100000001011" => data <= "000000";
				when "000100100000001100" => data <= "000000";
				when "000100100000001101" => data <= "000000";
				when "000100100000001110" => data <= "000000";
				when "000100100000001111" => data <= "000000";
				when "000100100000010000" => data <= "000000";
				when "000100100000010001" => data <= "000000";
				when "000100100000010010" => data <= "000000";
				when "000100100000010011" => data <= "000000";
				when "000100100000010100" => data <= "000000";
				when "000100100000010101" => data <= "000000";
				when "000100100000010110" => data <= "000000";
				when "000100100000010111" => data <= "000000";
				when "000100100000011000" => data <= "000000";
				when "000100100000011001" => data <= "000000";
				when "000100100000011010" => data <= "000000";
				when "000100100000011011" => data <= "000000";
				when "000100100000011100" => data <= "000000";
				when "000100100000011101" => data <= "000000";
				when "000100100000011110" => data <= "000000";
				when "000100100000011111" => data <= "000000";
				when "000100100000100000" => data <= "000000";
				when "000100100000100001" => data <= "000000";
				when "000100100000100010" => data <= "000000";
				when "000100100000100011" => data <= "000000";
				when "000100100000100100" => data <= "000000";
				when "000100100000100101" => data <= "000000";
				when "000100100000100110" => data <= "000000";
				when "000100100000100111" => data <= "000000";
				when "000100100000101000" => data <= "000000";
				when "000100100000101001" => data <= "000000";
				when "000100100000101010" => data <= "000000";
				when "000100100000101011" => data <= "000000";
				when "000100100000101100" => data <= "000000";
				when "000100100000101101" => data <= "000000";
				when "000100100000101110" => data <= "000000";
				when "000100100000101111" => data <= "000000";
				when "000100100000110000" => data <= "000000";
				when "000100100000110001" => data <= "000000";
				when "000100100000110010" => data <= "000000";
				when "000100100000110011" => data <= "000000";
				when "000100100000110100" => data <= "000000";
				when "000100100000110101" => data <= "000000";
				when "000100100000110110" => data <= "000000";
				when "000100100000110111" => data <= "000000";
				when "000100100000111000" => data <= "000000";
				when "000100100000111001" => data <= "000000";
				when "000100100000111010" => data <= "000000";
				when "000100100000111011" => data <= "000000";
				when "000100100000111100" => data <= "000000";
				when "000100100000111101" => data <= "000000";
				when "000100100000111110" => data <= "000000";
				when "000100100000111111" => data <= "000000";
				when "000100100001000000" => data <= "000000";
				when "000100100001000001" => data <= "000000";
				when "000100100001000010" => data <= "000000";
				when "000100100001000011" => data <= "000000";
				when "000100100001000100" => data <= "000000";
				when "000100100001000101" => data <= "000000";
				when "000100100001000110" => data <= "000000";
				when "000100100001000111" => data <= "000000";
				when "000100100001001000" => data <= "000000";
				when "000100100001001001" => data <= "000000";
				when "000100100001001010" => data <= "000000";
				when "000100100001001011" => data <= "000000";
				when "000100100001001100" => data <= "000000";
				when "000100100001001101" => data <= "000000";
				when "000100100001001110" => data <= "000000";
				when "000100100001001111" => data <= "000000";
				when "000100100001010000" => data <= "000000";
				when "000100100001010001" => data <= "000000";
				when "000100100001010010" => data <= "000000";
				when "000100100001010011" => data <= "000000";
				when "000100100001010100" => data <= "000000";
				when "000100100001010101" => data <= "000000";
				when "000100100001010110" => data <= "000000";
				when "000100100001010111" => data <= "000000";
				when "000100100001011000" => data <= "000000";
				when "000100100001011001" => data <= "000000";
				when "000100100001011010" => data <= "000000";
				when "000100100001011011" => data <= "000000";
				when "000100100001011100" => data <= "000000";
				when "000100100001011101" => data <= "000000";
				when "000100100001011110" => data <= "000000";
				when "000100100001011111" => data <= "000000";
				when "000100100001100000" => data <= "000000";
				when "000100100001100001" => data <= "000000";
				when "000100100001100010" => data <= "000000";
				when "000100100001100011" => data <= "000000";
				when "000100100001100100" => data <= "000000";
				when "000100100001100101" => data <= "000000";
				when "000100100001100110" => data <= "000000";
				when "000100100001100111" => data <= "000000";
				when "000100100001101000" => data <= "000000";
				when "000100100001101001" => data <= "000000";
				when "000100100001101010" => data <= "000000";
				when "000100100001101011" => data <= "000000";
				when "000100100001101100" => data <= "000000";
				when "000100100001101101" => data <= "000000";
				when "000100100001101110" => data <= "000000";
				when "000100100001101111" => data <= "000000";
				when "000100100001110000" => data <= "000000";
				when "000100100001110001" => data <= "000000";
				when "000100100001110010" => data <= "000000";
				when "000100100001110011" => data <= "000000";
				when "000100100001110100" => data <= "000000";
				when "000100100001110101" => data <= "000000";
				when "000100100001110110" => data <= "000000";
				when "000100100001110111" => data <= "000000";
				when "000100100001111000" => data <= "000000";
				when "000100100001111001" => data <= "000000";
				when "000100100001111010" => data <= "000000";
				when "000100100001111011" => data <= "000000";
				when "000100100001111100" => data <= "000000";
				when "000100100001111101" => data <= "000000";
				when "000100100001111110" => data <= "000000";
				when "000100100001111111" => data <= "000000";
				when "000100100010000000" => data <= "000000";
				when "000100100010000001" => data <= "000000";
				when "000100100010000010" => data <= "000000";
				when "000100100010000011" => data <= "000000";
				when "000100100010000100" => data <= "000000";
				when "000100100010000101" => data <= "000000";
				when "000100100010000110" => data <= "000000";
				when "000100100010000111" => data <= "000000";
				when "000100100010001000" => data <= "000000";
				when "000100100010001001" => data <= "000000";
				when "000100100010001010" => data <= "000000";
				when "000100100010001011" => data <= "000000";
				when "000100100010001100" => data <= "000000";
				when "000100100010001101" => data <= "000000";
				when "000100100010001110" => data <= "000000";
				when "000100100010001111" => data <= "000000";
				when "000100100010010000" => data <= "000000";
				when "000100100010010001" => data <= "000000";
				when "000100100010010010" => data <= "000000";
				when "000100100010010011" => data <= "000000";
				when "000100100010010100" => data <= "000000";
				when "000100100010010101" => data <= "000000";
				when "000100100010010110" => data <= "000000";
				when "000100100010010111" => data <= "000000";
				when "000100100010011000" => data <= "000000";
				when "000100100010011001" => data <= "000000";
				when "000100100010011010" => data <= "000000";
				when "000100100010011011" => data <= "000000";
				when "000100100010011100" => data <= "000000";
				when "000100100010011101" => data <= "000000";
				when "000100100010011110" => data <= "000000";
				when "000100100010011111" => data <= "000000";
				when "000100101000000000" => data <= "000000";
				when "000100101000000001" => data <= "000000";
				when "000100101000000010" => data <= "000000";
				when "000100101000000011" => data <= "000000";
				when "000100101000000100" => data <= "000000";
				when "000100101000000101" => data <= "000000";
				when "000100101000000110" => data <= "000000";
				when "000100101000000111" => data <= "000000";
				when "000100101000001000" => data <= "000000";
				when "000100101000001001" => data <= "000000";
				when "000100101000001010" => data <= "000000";
				when "000100101000001011" => data <= "000000";
				when "000100101000001100" => data <= "000000";
				when "000100101000001101" => data <= "000000";
				when "000100101000001110" => data <= "000000";
				when "000100101000001111" => data <= "000000";
				when "000100101000010000" => data <= "000000";
				when "000100101000010001" => data <= "000000";
				when "000100101000010010" => data <= "000000";
				when "000100101000010011" => data <= "000000";
				when "000100101000010100" => data <= "000000";
				when "000100101000010101" => data <= "000000";
				when "000100101000010110" => data <= "000000";
				when "000100101000010111" => data <= "000000";
				when "000100101000011000" => data <= "000000";
				when "000100101000011001" => data <= "000000";
				when "000100101000011010" => data <= "000000";
				when "000100101000011011" => data <= "000000";
				when "000100101000011100" => data <= "000000";
				when "000100101000011101" => data <= "000000";
				when "000100101000011110" => data <= "000000";
				when "000100101000011111" => data <= "000000";
				when "000100101000100000" => data <= "000000";
				when "000100101000100001" => data <= "000000";
				when "000100101000100010" => data <= "000000";
				when "000100101000100011" => data <= "000000";
				when "000100101000100100" => data <= "000000";
				when "000100101000100101" => data <= "000000";
				when "000100101000100110" => data <= "000000";
				when "000100101000100111" => data <= "000000";
				when "000100101000101000" => data <= "000000";
				when "000100101000101001" => data <= "000000";
				when "000100101000101010" => data <= "000000";
				when "000100101000101011" => data <= "000000";
				when "000100101000101100" => data <= "000000";
				when "000100101000101101" => data <= "000000";
				when "000100101000101110" => data <= "000000";
				when "000100101000101111" => data <= "000000";
				when "000100101000110000" => data <= "000000";
				when "000100101000110001" => data <= "000000";
				when "000100101000110010" => data <= "000000";
				when "000100101000110011" => data <= "000000";
				when "000100101000110100" => data <= "000000";
				when "000100101000110101" => data <= "000000";
				when "000100101000110110" => data <= "000000";
				when "000100101000110111" => data <= "000000";
				when "000100101000111000" => data <= "000000";
				when "000100101000111001" => data <= "000000";
				when "000100101000111010" => data <= "000000";
				when "000100101000111011" => data <= "000000";
				when "000100101000111100" => data <= "000000";
				when "000100101000111101" => data <= "000000";
				when "000100101000111110" => data <= "000000";
				when "000100101000111111" => data <= "000000";
				when "000100101001000000" => data <= "000000";
				when "000100101001000001" => data <= "000000";
				when "000100101001000010" => data <= "000000";
				when "000100101001000011" => data <= "000000";
				when "000100101001000100" => data <= "000000";
				when "000100101001000101" => data <= "000000";
				when "000100101001000110" => data <= "000000";
				when "000100101001000111" => data <= "000000";
				when "000100101001001000" => data <= "000000";
				when "000100101001001001" => data <= "000000";
				when "000100101001001010" => data <= "000000";
				when "000100101001001011" => data <= "000000";
				when "000100101001001100" => data <= "000000";
				when "000100101001001101" => data <= "000000";
				when "000100101001001110" => data <= "000000";
				when "000100101001001111" => data <= "000000";
				when "000100101001010000" => data <= "000000";
				when "000100101001010001" => data <= "000000";
				when "000100101001010010" => data <= "000000";
				when "000100101001010011" => data <= "000000";
				when "000100101001010100" => data <= "000000";
				when "000100101001010101" => data <= "000000";
				when "000100101001010110" => data <= "000000";
				when "000100101001010111" => data <= "000000";
				when "000100101001011000" => data <= "000000";
				when "000100101001011001" => data <= "000000";
				when "000100101001011010" => data <= "000000";
				when "000100101001011011" => data <= "000000";
				when "000100101001011100" => data <= "000000";
				when "000100101001011101" => data <= "000000";
				when "000100101001011110" => data <= "000000";
				when "000100101001011111" => data <= "000000";
				when "000100101001100000" => data <= "000000";
				when "000100101001100001" => data <= "000000";
				when "000100101001100010" => data <= "000000";
				when "000100101001100011" => data <= "000000";
				when "000100101001100100" => data <= "000000";
				when "000100101001100101" => data <= "000000";
				when "000100101001100110" => data <= "000000";
				when "000100101001100111" => data <= "000000";
				when "000100101001101000" => data <= "000000";
				when "000100101001101001" => data <= "000000";
				when "000100101001101010" => data <= "000000";
				when "000100101001101011" => data <= "000000";
				when "000100101001101100" => data <= "000000";
				when "000100101001101101" => data <= "000000";
				when "000100101001101110" => data <= "000000";
				when "000100101001101111" => data <= "000000";
				when "000100101001110000" => data <= "000000";
				when "000100101001110001" => data <= "000000";
				when "000100101001110010" => data <= "000000";
				when "000100101001110011" => data <= "000000";
				when "000100101001110100" => data <= "000000";
				when "000100101001110101" => data <= "000000";
				when "000100101001110110" => data <= "000000";
				when "000100101001110111" => data <= "000000";
				when "000100101001111000" => data <= "000000";
				when "000100101001111001" => data <= "000000";
				when "000100101001111010" => data <= "000000";
				when "000100101001111011" => data <= "000000";
				when "000100101001111100" => data <= "000000";
				when "000100101001111101" => data <= "000000";
				when "000100101001111110" => data <= "000000";
				when "000100101001111111" => data <= "000000";
				when "000100101010000000" => data <= "000000";
				when "000100101010000001" => data <= "000000";
				when "000100101010000010" => data <= "000000";
				when "000100101010000011" => data <= "000000";
				when "000100101010000100" => data <= "000000";
				when "000100101010000101" => data <= "000000";
				when "000100101010000110" => data <= "000000";
				when "000100101010000111" => data <= "000000";
				when "000100101010001000" => data <= "000000";
				when "000100101010001001" => data <= "000000";
				when "000100101010001010" => data <= "000000";
				when "000100101010001011" => data <= "000000";
				when "000100101010001100" => data <= "000000";
				when "000100101010001101" => data <= "000000";
				when "000100101010001110" => data <= "000000";
				when "000100101010001111" => data <= "000000";
				when "000100101010010000" => data <= "000000";
				when "000100101010010001" => data <= "000000";
				when "000100101010010010" => data <= "000000";
				when "000100101010010011" => data <= "000000";
				when "000100101010010100" => data <= "000000";
				when "000100101010010101" => data <= "000000";
				when "000100101010010110" => data <= "000000";
				when "000100101010010111" => data <= "000000";
				when "000100101010011000" => data <= "000000";
				when "000100101010011001" => data <= "000000";
				when "000100101010011010" => data <= "000000";
				when "000100101010011011" => data <= "000000";
				when "000100101010011100" => data <= "000000";
				when "000100101010011101" => data <= "000000";
				when "000100101010011110" => data <= "000000";
				when "000100101010011111" => data <= "000000";
				when "000100110000000000" => data <= "000000";
				when "000100110000000001" => data <= "000000";
				when "000100110000000010" => data <= "000000";
				when "000100110000000011" => data <= "000000";
				when "000100110000000100" => data <= "000000";
				when "000100110000000101" => data <= "000000";
				when "000100110000000110" => data <= "000000";
				when "000100110000000111" => data <= "000000";
				when "000100110000001000" => data <= "000000";
				when "000100110000001001" => data <= "000000";
				when "000100110000001010" => data <= "000000";
				when "000100110000001011" => data <= "000000";
				when "000100110000001100" => data <= "000000";
				when "000100110000001101" => data <= "000000";
				when "000100110000001110" => data <= "000000";
				when "000100110000001111" => data <= "000000";
				when "000100110000010000" => data <= "000000";
				when "000100110000010001" => data <= "000000";
				when "000100110000010010" => data <= "000000";
				when "000100110000010011" => data <= "000000";
				when "000100110000010100" => data <= "000000";
				when "000100110000010101" => data <= "000000";
				when "000100110000010110" => data <= "000000";
				when "000100110000010111" => data <= "000000";
				when "000100110000011000" => data <= "000000";
				when "000100110000011001" => data <= "000000";
				when "000100110000011010" => data <= "000000";
				when "000100110000011011" => data <= "000000";
				when "000100110000011100" => data <= "000000";
				when "000100110000011101" => data <= "000000";
				when "000100110000011110" => data <= "000000";
				when "000100110000011111" => data <= "000000";
				when "000100110000100000" => data <= "000000";
				when "000100110000100001" => data <= "000000";
				when "000100110000100010" => data <= "000000";
				when "000100110000100011" => data <= "000000";
				when "000100110000100100" => data <= "000000";
				when "000100110000100101" => data <= "000000";
				when "000100110000100110" => data <= "000000";
				when "000100110000100111" => data <= "000000";
				when "000100110000101000" => data <= "000000";
				when "000100110000101001" => data <= "000000";
				when "000100110000101010" => data <= "000000";
				when "000100110000101011" => data <= "000000";
				when "000100110000101100" => data <= "000000";
				when "000100110000101101" => data <= "000000";
				when "000100110000101110" => data <= "000000";
				when "000100110000101111" => data <= "000000";
				when "000100110000110000" => data <= "000000";
				when "000100110000110001" => data <= "000000";
				when "000100110000110010" => data <= "000000";
				when "000100110000110011" => data <= "000000";
				when "000100110000110100" => data <= "000000";
				when "000100110000110101" => data <= "000000";
				when "000100110000110110" => data <= "000000";
				when "000100110000110111" => data <= "000000";
				when "000100110000111000" => data <= "000000";
				when "000100110000111001" => data <= "000000";
				when "000100110000111010" => data <= "000000";
				when "000100110000111011" => data <= "000000";
				when "000100110000111100" => data <= "000000";
				when "000100110000111101" => data <= "000000";
				when "000100110000111110" => data <= "000000";
				when "000100110000111111" => data <= "000000";
				when "000100110001000000" => data <= "000000";
				when "000100110001000001" => data <= "000000";
				when "000100110001000010" => data <= "000000";
				when "000100110001000011" => data <= "000000";
				when "000100110001000100" => data <= "000000";
				when "000100110001000101" => data <= "000000";
				when "000100110001000110" => data <= "000000";
				when "000100110001000111" => data <= "000000";
				when "000100110001001000" => data <= "000000";
				when "000100110001001001" => data <= "000000";
				when "000100110001001010" => data <= "000000";
				when "000100110001001011" => data <= "000000";
				when "000100110001001100" => data <= "000000";
				when "000100110001001101" => data <= "000000";
				when "000100110001001110" => data <= "000000";
				when "000100110001001111" => data <= "000000";
				when "000100110001010000" => data <= "000000";
				when "000100110001010001" => data <= "000000";
				when "000100110001010010" => data <= "000000";
				when "000100110001010011" => data <= "000000";
				when "000100110001010100" => data <= "000000";
				when "000100110001010101" => data <= "000000";
				when "000100110001010110" => data <= "000000";
				when "000100110001010111" => data <= "000000";
				when "000100110001011000" => data <= "000000";
				when "000100110001011001" => data <= "000000";
				when "000100110001011010" => data <= "000000";
				when "000100110001011011" => data <= "000000";
				when "000100110001011100" => data <= "000000";
				when "000100110001011101" => data <= "000000";
				when "000100110001011110" => data <= "000000";
				when "000100110001011111" => data <= "000000";
				when "000100110001100000" => data <= "000000";
				when "000100110001100001" => data <= "000000";
				when "000100110001100010" => data <= "000000";
				when "000100110001100011" => data <= "000000";
				when "000100110001100100" => data <= "000000";
				when "000100110001100101" => data <= "000000";
				when "000100110001100110" => data <= "000000";
				when "000100110001100111" => data <= "000000";
				when "000100110001101000" => data <= "000000";
				when "000100110001101001" => data <= "000000";
				when "000100110001101010" => data <= "000000";
				when "000100110001101011" => data <= "000000";
				when "000100110001101100" => data <= "000000";
				when "000100110001101101" => data <= "000000";
				when "000100110001101110" => data <= "000000";
				when "000100110001101111" => data <= "000000";
				when "000100110001110000" => data <= "000000";
				when "000100110001110001" => data <= "000000";
				when "000100110001110010" => data <= "000000";
				when "000100110001110011" => data <= "000000";
				when "000100110001110100" => data <= "000000";
				when "000100110001110101" => data <= "000000";
				when "000100110001110110" => data <= "000000";
				when "000100110001110111" => data <= "000000";
				when "000100110001111000" => data <= "000000";
				when "000100110001111001" => data <= "000000";
				when "000100110001111010" => data <= "000000";
				when "000100110001111011" => data <= "000000";
				when "000100110001111100" => data <= "000000";
				when "000100110001111101" => data <= "000000";
				when "000100110001111110" => data <= "000000";
				when "000100110001111111" => data <= "000000";
				when "000100110010000000" => data <= "000000";
				when "000100110010000001" => data <= "000000";
				when "000100110010000010" => data <= "000000";
				when "000100110010000011" => data <= "000000";
				when "000100110010000100" => data <= "000000";
				when "000100110010000101" => data <= "000000";
				when "000100110010000110" => data <= "000000";
				when "000100110010000111" => data <= "000000";
				when "000100110010001000" => data <= "000000";
				when "000100110010001001" => data <= "000000";
				when "000100110010001010" => data <= "000000";
				when "000100110010001011" => data <= "000000";
				when "000100110010001100" => data <= "000000";
				when "000100110010001101" => data <= "000000";
				when "000100110010001110" => data <= "000000";
				when "000100110010001111" => data <= "000000";
				when "000100110010010000" => data <= "000000";
				when "000100110010010001" => data <= "000000";
				when "000100110010010010" => data <= "000000";
				when "000100110010010011" => data <= "000000";
				when "000100110010010100" => data <= "000000";
				when "000100110010010101" => data <= "000000";
				when "000100110010010110" => data <= "000000";
				when "000100110010010111" => data <= "000000";
				when "000100110010011000" => data <= "000000";
				when "000100110010011001" => data <= "000000";
				when "000100110010011010" => data <= "000000";
				when "000100110010011011" => data <= "000000";
				when "000100110010011100" => data <= "000000";
				when "000100110010011101" => data <= "000000";
				when "000100110010011110" => data <= "000000";
				when "000100110010011111" => data <= "000000";
				when "000100111000000000" => data <= "000000";
				when "000100111000000001" => data <= "000000";
				when "000100111000000010" => data <= "000000";
				when "000100111000000011" => data <= "000000";
				when "000100111000000100" => data <= "000000";
				when "000100111000000101" => data <= "000000";
				when "000100111000000110" => data <= "000000";
				when "000100111000000111" => data <= "000000";
				when "000100111000001000" => data <= "000000";
				when "000100111000001001" => data <= "000000";
				when "000100111000001010" => data <= "000000";
				when "000100111000001011" => data <= "000000";
				when "000100111000001100" => data <= "000000";
				when "000100111000001101" => data <= "000000";
				when "000100111000001110" => data <= "000000";
				when "000100111000001111" => data <= "000000";
				when "000100111000010000" => data <= "000000";
				when "000100111000010001" => data <= "000000";
				when "000100111000010010" => data <= "000000";
				when "000100111000010011" => data <= "000000";
				when "000100111000010100" => data <= "000000";
				when "000100111000010101" => data <= "000000";
				when "000100111000010110" => data <= "000000";
				when "000100111000010111" => data <= "000000";
				when "000100111000011000" => data <= "000000";
				when "000100111000011001" => data <= "000000";
				when "000100111000011010" => data <= "000000";
				when "000100111000011011" => data <= "000000";
				when "000100111000011100" => data <= "000000";
				when "000100111000011101" => data <= "000000";
				when "000100111000011110" => data <= "000000";
				when "000100111000011111" => data <= "000000";
				when "000100111000100000" => data <= "000000";
				when "000100111000100001" => data <= "000000";
				when "000100111000100010" => data <= "000000";
				when "000100111000100011" => data <= "000000";
				when "000100111000100100" => data <= "000000";
				when "000100111000100101" => data <= "000000";
				when "000100111000100110" => data <= "000000";
				when "000100111000100111" => data <= "000000";
				when "000100111000101000" => data <= "000000";
				when "000100111000101001" => data <= "000000";
				when "000100111000101010" => data <= "000000";
				when "000100111000101011" => data <= "000000";
				when "000100111000101100" => data <= "000000";
				when "000100111000101101" => data <= "000000";
				when "000100111000101110" => data <= "000000";
				when "000100111000101111" => data <= "000000";
				when "000100111000110000" => data <= "000000";
				when "000100111000110001" => data <= "000000";
				when "000100111000110010" => data <= "000000";
				when "000100111000110011" => data <= "000000";
				when "000100111000110100" => data <= "000000";
				when "000100111000110101" => data <= "000000";
				when "000100111000110110" => data <= "000000";
				when "000100111000110111" => data <= "000000";
				when "000100111000111000" => data <= "000000";
				when "000100111000111001" => data <= "000000";
				when "000100111000111010" => data <= "000000";
				when "000100111000111011" => data <= "000000";
				when "000100111000111100" => data <= "000000";
				when "000100111000111101" => data <= "000000";
				when "000100111000111110" => data <= "000000";
				when "000100111000111111" => data <= "000000";
				when "000100111001000000" => data <= "000000";
				when "000100111001000001" => data <= "000000";
				when "000100111001000010" => data <= "000000";
				when "000100111001000011" => data <= "000000";
				when "000100111001000100" => data <= "000000";
				when "000100111001000101" => data <= "000000";
				when "000100111001000110" => data <= "000000";
				when "000100111001000111" => data <= "000000";
				when "000100111001001000" => data <= "000000";
				when "000100111001001001" => data <= "000000";
				when "000100111001001010" => data <= "000000";
				when "000100111001001011" => data <= "000000";
				when "000100111001001100" => data <= "000000";
				when "000100111001001101" => data <= "000000";
				when "000100111001001110" => data <= "000000";
				when "000100111001001111" => data <= "000000";
				when "000100111001010000" => data <= "000000";
				when "000100111001010001" => data <= "000000";
				when "000100111001010010" => data <= "000000";
				when "000100111001010011" => data <= "000000";
				when "000100111001010100" => data <= "000000";
				when "000100111001010101" => data <= "000000";
				when "000100111001010110" => data <= "000000";
				when "000100111001010111" => data <= "000000";
				when "000100111001011000" => data <= "000000";
				when "000100111001011001" => data <= "000000";
				when "000100111001011010" => data <= "000000";
				when "000100111001011011" => data <= "000000";
				when "000100111001011100" => data <= "000000";
				when "000100111001011101" => data <= "000000";
				when "000100111001011110" => data <= "000000";
				when "000100111001011111" => data <= "000000";
				when "000100111001100000" => data <= "000000";
				when "000100111001100001" => data <= "000000";
				when "000100111001100010" => data <= "000000";
				when "000100111001100011" => data <= "000000";
				when "000100111001100100" => data <= "000000";
				when "000100111001100101" => data <= "000000";
				when "000100111001100110" => data <= "000000";
				when "000100111001100111" => data <= "000000";
				when "000100111001101000" => data <= "000000";
				when "000100111001101001" => data <= "000000";
				when "000100111001101010" => data <= "000000";
				when "000100111001101011" => data <= "000000";
				when "000100111001101100" => data <= "000000";
				when "000100111001101101" => data <= "000000";
				when "000100111001101110" => data <= "000000";
				when "000100111001101111" => data <= "000000";
				when "000100111001110000" => data <= "000000";
				when "000100111001110001" => data <= "000000";
				when "000100111001110010" => data <= "000000";
				when "000100111001110011" => data <= "000000";
				when "000100111001110100" => data <= "000000";
				when "000100111001110101" => data <= "000000";
				when "000100111001110110" => data <= "000000";
				when "000100111001110111" => data <= "000000";
				when "000100111001111000" => data <= "000000";
				when "000100111001111001" => data <= "000000";
				when "000100111001111010" => data <= "000000";
				when "000100111001111011" => data <= "000000";
				when "000100111001111100" => data <= "000000";
				when "000100111001111101" => data <= "000000";
				when "000100111001111110" => data <= "000000";
				when "000100111001111111" => data <= "000000";
				when "000100111010000000" => data <= "000000";
				when "000100111010000001" => data <= "000000";
				when "000100111010000010" => data <= "000000";
				when "000100111010000011" => data <= "000000";
				when "000100111010000100" => data <= "000000";
				when "000100111010000101" => data <= "000000";
				when "000100111010000110" => data <= "000000";
				when "000100111010000111" => data <= "000000";
				when "000100111010001000" => data <= "000000";
				when "000100111010001001" => data <= "000000";
				when "000100111010001010" => data <= "000000";
				when "000100111010001011" => data <= "000000";
				when "000100111010001100" => data <= "000000";
				when "000100111010001101" => data <= "000000";
				when "000100111010001110" => data <= "000000";
				when "000100111010001111" => data <= "000000";
				when "000100111010010000" => data <= "000000";
				when "000100111010010001" => data <= "000000";
				when "000100111010010010" => data <= "000000";
				when "000100111010010011" => data <= "000000";
				when "000100111010010100" => data <= "000000";
				when "000100111010010101" => data <= "000000";
				when "000100111010010110" => data <= "000000";
				when "000100111010010111" => data <= "000000";
				when "000100111010011000" => data <= "000000";
				when "000100111010011001" => data <= "000000";
				when "000100111010011010" => data <= "000000";
				when "000100111010011011" => data <= "000000";
				when "000100111010011100" => data <= "000000";
				when "000100111010011101" => data <= "000000";
				when "000100111010011110" => data <= "000000";
				when "000100111010011111" => data <= "000000";
				when "000101000000000000" => data <= "000000";
				when "000101000000000001" => data <= "000000";
				when "000101000000000010" => data <= "000000";
				when "000101000000000011" => data <= "000000";
				when "000101000000000100" => data <= "000000";
				when "000101000000000101" => data <= "000000";
				when "000101000000000110" => data <= "000000";
				when "000101000000000111" => data <= "000000";
				when "000101000000001000" => data <= "000000";
				when "000101000000001001" => data <= "000000";
				when "000101000000001010" => data <= "000000";
				when "000101000000001011" => data <= "000000";
				when "000101000000001100" => data <= "000000";
				when "000101000000001101" => data <= "000000";
				when "000101000000001110" => data <= "000000";
				when "000101000000001111" => data <= "000000";
				when "000101000000010000" => data <= "000000";
				when "000101000000010001" => data <= "000000";
				when "000101000000010010" => data <= "000000";
				when "000101000000010011" => data <= "000000";
				when "000101000000010100" => data <= "000000";
				when "000101000000010101" => data <= "000000";
				when "000101000000010110" => data <= "000000";
				when "000101000000010111" => data <= "000000";
				when "000101000000011000" => data <= "000000";
				when "000101000000011001" => data <= "000000";
				when "000101000000011010" => data <= "000000";
				when "000101000000011011" => data <= "000000";
				when "000101000000011100" => data <= "000000";
				when "000101000000011101" => data <= "000000";
				when "000101000000011110" => data <= "000000";
				when "000101000000011111" => data <= "000000";
				when "000101000000100000" => data <= "000000";
				when "000101000000100001" => data <= "000000";
				when "000101000000100010" => data <= "000000";
				when "000101000000100011" => data <= "000000";
				when "000101000000100100" => data <= "000000";
				when "000101000000100101" => data <= "000000";
				when "000101000000100110" => data <= "000000";
				when "000101000000100111" => data <= "000000";
				when "000101000000101000" => data <= "000000";
				when "000101000000101001" => data <= "000000";
				when "000101000000101010" => data <= "000000";
				when "000101000000101011" => data <= "000000";
				when "000101000000101100" => data <= "000000";
				when "000101000000101101" => data <= "000000";
				when "000101000000101110" => data <= "000000";
				when "000101000000101111" => data <= "000000";
				when "000101000000110000" => data <= "000000";
				when "000101000000110001" => data <= "000000";
				when "000101000000110010" => data <= "000000";
				when "000101000000110011" => data <= "000000";
				when "000101000000110100" => data <= "000000";
				when "000101000000110101" => data <= "000000";
				when "000101000000110110" => data <= "000000";
				when "000101000000110111" => data <= "000000";
				when "000101000000111000" => data <= "000000";
				when "000101000000111001" => data <= "000000";
				when "000101000000111010" => data <= "000000";
				when "000101000000111011" => data <= "000000";
				when "000101000000111100" => data <= "000000";
				when "000101000000111101" => data <= "000000";
				when "000101000000111110" => data <= "000000";
				when "000101000000111111" => data <= "000000";
				when "000101000001000000" => data <= "000000";
				when "000101000001000001" => data <= "000000";
				when "000101000001000010" => data <= "000000";
				when "000101000001000011" => data <= "000000";
				when "000101000001000100" => data <= "000000";
				when "000101000001000101" => data <= "000000";
				when "000101000001000110" => data <= "000000";
				when "000101000001000111" => data <= "000000";
				when "000101000001001000" => data <= "000000";
				when "000101000001001001" => data <= "000000";
				when "000101000001001010" => data <= "000000";
				when "000101000001001011" => data <= "000000";
				when "000101000001001100" => data <= "000000";
				when "000101000001001101" => data <= "000000";
				when "000101000001001110" => data <= "000000";
				when "000101000001001111" => data <= "000000";
				when "000101000001010000" => data <= "000000";
				when "000101000001010001" => data <= "000000";
				when "000101000001010010" => data <= "000000";
				when "000101000001010011" => data <= "000000";
				when "000101000001010100" => data <= "000000";
				when "000101000001010101" => data <= "000000";
				when "000101000001010110" => data <= "000000";
				when "000101000001010111" => data <= "000000";
				when "000101000001011000" => data <= "000000";
				when "000101000001011001" => data <= "000000";
				when "000101000001011010" => data <= "000000";
				when "000101000001011011" => data <= "000000";
				when "000101000001011100" => data <= "000000";
				when "000101000001011101" => data <= "000000";
				when "000101000001011110" => data <= "000000";
				when "000101000001011111" => data <= "000000";
				when "000101000001100000" => data <= "000000";
				when "000101000001100001" => data <= "000000";
				when "000101000001100010" => data <= "000000";
				when "000101000001100011" => data <= "000000";
				when "000101000001100100" => data <= "000000";
				when "000101000001100101" => data <= "000000";
				when "000101000001100110" => data <= "000000";
				when "000101000001100111" => data <= "000000";
				when "000101000001101000" => data <= "000000";
				when "000101000001101001" => data <= "000000";
				when "000101000001101010" => data <= "000000";
				when "000101000001101011" => data <= "000000";
				when "000101000001101100" => data <= "000000";
				when "000101000001101101" => data <= "000000";
				when "000101000001101110" => data <= "000000";
				when "000101000001101111" => data <= "000000";
				when "000101000001110000" => data <= "000000";
				when "000101000001110001" => data <= "000000";
				when "000101000001110010" => data <= "000000";
				when "000101000001110011" => data <= "000000";
				when "000101000001110100" => data <= "000000";
				when "000101000001110101" => data <= "000000";
				when "000101000001110110" => data <= "000000";
				when "000101000001110111" => data <= "000000";
				when "000101000001111000" => data <= "000000";
				when "000101000001111001" => data <= "000000";
				when "000101000001111010" => data <= "000000";
				when "000101000001111011" => data <= "000000";
				when "000101000001111100" => data <= "000000";
				when "000101000001111101" => data <= "000000";
				when "000101000001111110" => data <= "000000";
				when "000101000001111111" => data <= "000000";
				when "000101000010000000" => data <= "000000";
				when "000101000010000001" => data <= "000000";
				when "000101000010000010" => data <= "000000";
				when "000101000010000011" => data <= "000000";
				when "000101000010000100" => data <= "000000";
				when "000101000010000101" => data <= "000000";
				when "000101000010000110" => data <= "000000";
				when "000101000010000111" => data <= "000000";
				when "000101000010001000" => data <= "000000";
				when "000101000010001001" => data <= "000000";
				when "000101000010001010" => data <= "000000";
				when "000101000010001011" => data <= "000000";
				when "000101000010001100" => data <= "000000";
				when "000101000010001101" => data <= "000000";
				when "000101000010001110" => data <= "000000";
				when "000101000010001111" => data <= "000000";
				when "000101000010010000" => data <= "000000";
				when "000101000010010001" => data <= "000000";
				when "000101000010010010" => data <= "000000";
				when "000101000010010011" => data <= "000000";
				when "000101000010010100" => data <= "000000";
				when "000101000010010101" => data <= "000000";
				when "000101000010010110" => data <= "000000";
				when "000101000010010111" => data <= "000000";
				when "000101000010011000" => data <= "000000";
				when "000101000010011001" => data <= "000000";
				when "000101000010011010" => data <= "000000";
				when "000101000010011011" => data <= "000000";
				when "000101000010011100" => data <= "000000";
				when "000101000010011101" => data <= "000000";
				when "000101000010011110" => data <= "000000";
				when "000101000010011111" => data <= "000000";
				when "000101001000000000" => data <= "000000";
				when "000101001000000001" => data <= "000000";
				when "000101001000000010" => data <= "000000";
				when "000101001000000011" => data <= "000000";
				when "000101001000000100" => data <= "000000";
				when "000101001000000101" => data <= "000000";
				when "000101001000000110" => data <= "000000";
				when "000101001000000111" => data <= "000000";
				when "000101001000001000" => data <= "000000";
				when "000101001000001001" => data <= "000000";
				when "000101001000001010" => data <= "000000";
				when "000101001000001011" => data <= "000000";
				when "000101001000001100" => data <= "000000";
				when "000101001000001101" => data <= "000000";
				when "000101001000001110" => data <= "000000";
				when "000101001000001111" => data <= "000000";
				when "000101001000010000" => data <= "000000";
				when "000101001000010001" => data <= "000000";
				when "000101001000010010" => data <= "000000";
				when "000101001000010011" => data <= "000000";
				when "000101001000010100" => data <= "000000";
				when "000101001000010101" => data <= "000000";
				when "000101001000010110" => data <= "000000";
				when "000101001000010111" => data <= "000000";
				when "000101001000011000" => data <= "000000";
				when "000101001000011001" => data <= "000000";
				when "000101001000011010" => data <= "000000";
				when "000101001000011011" => data <= "000000";
				when "000101001000011100" => data <= "000000";
				when "000101001000011101" => data <= "000000";
				when "000101001000011110" => data <= "000000";
				when "000101001000011111" => data <= "000000";
				when "000101001000100000" => data <= "000000";
				when "000101001000100001" => data <= "000000";
				when "000101001000100010" => data <= "000000";
				when "000101001000100011" => data <= "000000";
				when "000101001000100100" => data <= "000000";
				when "000101001000100101" => data <= "000000";
				when "000101001000100110" => data <= "000000";
				when "000101001000100111" => data <= "000000";
				when "000101001000101000" => data <= "000000";
				when "000101001000101001" => data <= "000000";
				when "000101001000101010" => data <= "000000";
				when "000101001000101011" => data <= "000000";
				when "000101001000101100" => data <= "000000";
				when "000101001000101101" => data <= "000000";
				when "000101001000101110" => data <= "000000";
				when "000101001000101111" => data <= "000000";
				when "000101001000110000" => data <= "000000";
				when "000101001000110001" => data <= "000000";
				when "000101001000110010" => data <= "000000";
				when "000101001000110011" => data <= "000000";
				when "000101001000110100" => data <= "000000";
				when "000101001000110101" => data <= "000000";
				when "000101001000110110" => data <= "000000";
				when "000101001000110111" => data <= "000000";
				when "000101001000111000" => data <= "000000";
				when "000101001000111001" => data <= "000000";
				when "000101001000111010" => data <= "000000";
				when "000101001000111011" => data <= "000000";
				when "000101001000111100" => data <= "000000";
				when "000101001000111101" => data <= "000000";
				when "000101001000111110" => data <= "000000";
				when "000101001000111111" => data <= "000000";
				when "000101001001000000" => data <= "000000";
				when "000101001001000001" => data <= "000000";
				when "000101001001000010" => data <= "000000";
				when "000101001001000011" => data <= "000000";
				when "000101001001000100" => data <= "000000";
				when "000101001001000101" => data <= "000000";
				when "000101001001000110" => data <= "000000";
				when "000101001001000111" => data <= "000000";
				when "000101001001001000" => data <= "000000";
				when "000101001001001001" => data <= "000000";
				when "000101001001001010" => data <= "000000";
				when "000101001001001011" => data <= "000000";
				when "000101001001001100" => data <= "000000";
				when "000101001001001101" => data <= "000000";
				when "000101001001001110" => data <= "000000";
				when "000101001001001111" => data <= "000000";
				when "000101001001010000" => data <= "000000";
				when "000101001001010001" => data <= "000000";
				when "000101001001010010" => data <= "000000";
				when "000101001001010011" => data <= "000000";
				when "000101001001010100" => data <= "000000";
				when "000101001001010101" => data <= "000000";
				when "000101001001010110" => data <= "000000";
				when "000101001001010111" => data <= "000000";
				when "000101001001011000" => data <= "000000";
				when "000101001001011001" => data <= "000000";
				when "000101001001011010" => data <= "000000";
				when "000101001001011011" => data <= "000000";
				when "000101001001011100" => data <= "000000";
				when "000101001001011101" => data <= "000000";
				when "000101001001011110" => data <= "000000";
				when "000101001001011111" => data <= "000000";
				when "000101001001100000" => data <= "000000";
				when "000101001001100001" => data <= "000000";
				when "000101001001100010" => data <= "000000";
				when "000101001001100011" => data <= "000000";
				when "000101001001100100" => data <= "000000";
				when "000101001001100101" => data <= "000000";
				when "000101001001100110" => data <= "000000";
				when "000101001001100111" => data <= "000000";
				when "000101001001101000" => data <= "000000";
				when "000101001001101001" => data <= "000000";
				when "000101001001101010" => data <= "000000";
				when "000101001001101011" => data <= "000000";
				when "000101001001101100" => data <= "000000";
				when "000101001001101101" => data <= "000000";
				when "000101001001101110" => data <= "000000";
				when "000101001001101111" => data <= "000000";
				when "000101001001110000" => data <= "000000";
				when "000101001001110001" => data <= "000000";
				when "000101001001110010" => data <= "000000";
				when "000101001001110011" => data <= "000000";
				when "000101001001110100" => data <= "000000";
				when "000101001001110101" => data <= "000000";
				when "000101001001110110" => data <= "000000";
				when "000101001001110111" => data <= "000000";
				when "000101001001111000" => data <= "000000";
				when "000101001001111001" => data <= "000000";
				when "000101001001111010" => data <= "000000";
				when "000101001001111011" => data <= "000000";
				when "000101001001111100" => data <= "000000";
				when "000101001001111101" => data <= "000000";
				when "000101001001111110" => data <= "000000";
				when "000101001001111111" => data <= "000000";
				when "000101001010000000" => data <= "000000";
				when "000101001010000001" => data <= "000000";
				when "000101001010000010" => data <= "000000";
				when "000101001010000011" => data <= "000000";
				when "000101001010000100" => data <= "000000";
				when "000101001010000101" => data <= "000000";
				when "000101001010000110" => data <= "000000";
				when "000101001010000111" => data <= "000000";
				when "000101001010001000" => data <= "000000";
				when "000101001010001001" => data <= "000000";
				when "000101001010001010" => data <= "000000";
				when "000101001010001011" => data <= "000000";
				when "000101001010001100" => data <= "000000";
				when "000101001010001101" => data <= "000000";
				when "000101001010001110" => data <= "000000";
				when "000101001010001111" => data <= "000000";
				when "000101001010010000" => data <= "000000";
				when "000101001010010001" => data <= "000000";
				when "000101001010010010" => data <= "000000";
				when "000101001010010011" => data <= "000000";
				when "000101001010010100" => data <= "000000";
				when "000101001010010101" => data <= "000000";
				when "000101001010010110" => data <= "000000";
				when "000101001010010111" => data <= "000000";
				when "000101001010011000" => data <= "000000";
				when "000101001010011001" => data <= "000000";
				when "000101001010011010" => data <= "000000";
				when "000101001010011011" => data <= "000000";
				when "000101001010011100" => data <= "000000";
				when "000101001010011101" => data <= "000000";
				when "000101001010011110" => data <= "000000";
				when "000101001010011111" => data <= "000000";
				when "000101010000000000" => data <= "000000";
				when "000101010000000001" => data <= "000000";
				when "000101010000000010" => data <= "000000";
				when "000101010000000011" => data <= "000000";
				when "000101010000000100" => data <= "000000";
				when "000101010000000101" => data <= "000000";
				when "000101010000000110" => data <= "000000";
				when "000101010000000111" => data <= "000000";
				when "000101010000001000" => data <= "000000";
				when "000101010000001001" => data <= "000000";
				when "000101010000001010" => data <= "000000";
				when "000101010000001011" => data <= "000000";
				when "000101010000001100" => data <= "000000";
				when "000101010000001101" => data <= "000000";
				when "000101010000001110" => data <= "000000";
				when "000101010000001111" => data <= "000000";
				when "000101010000010000" => data <= "000000";
				when "000101010000010001" => data <= "000000";
				when "000101010000010010" => data <= "000000";
				when "000101010000010011" => data <= "000000";
				when "000101010000010100" => data <= "000000";
				when "000101010000010101" => data <= "000000";
				when "000101010000010110" => data <= "000000";
				when "000101010000010111" => data <= "000000";
				when "000101010000011000" => data <= "000000";
				when "000101010000011001" => data <= "000000";
				when "000101010000011010" => data <= "000000";
				when "000101010000011011" => data <= "000000";
				when "000101010000011100" => data <= "000000";
				when "000101010000011101" => data <= "000000";
				when "000101010000011110" => data <= "000000";
				when "000101010000011111" => data <= "000000";
				when "000101010000100000" => data <= "000000";
				when "000101010000100001" => data <= "000000";
				when "000101010000100010" => data <= "000000";
				when "000101010000100011" => data <= "000000";
				when "000101010000100100" => data <= "000000";
				when "000101010000100101" => data <= "000000";
				when "000101010000100110" => data <= "000000";
				when "000101010000100111" => data <= "000000";
				when "000101010000101000" => data <= "000000";
				when "000101010000101001" => data <= "000000";
				when "000101010000101010" => data <= "000000";
				when "000101010000101011" => data <= "000000";
				when "000101010000101100" => data <= "000000";
				when "000101010000101101" => data <= "000000";
				when "000101010000101110" => data <= "000000";
				when "000101010000101111" => data <= "000000";
				when "000101010000110000" => data <= "000000";
				when "000101010000110001" => data <= "000000";
				when "000101010000110010" => data <= "000000";
				when "000101010000110011" => data <= "000000";
				when "000101010000110100" => data <= "000000";
				when "000101010000110101" => data <= "000000";
				when "000101010000110110" => data <= "000000";
				when "000101010000110111" => data <= "000000";
				when "000101010000111000" => data <= "000000";
				when "000101010000111001" => data <= "000000";
				when "000101010000111010" => data <= "000000";
				when "000101010000111011" => data <= "000000";
				when "000101010000111100" => data <= "000000";
				when "000101010000111101" => data <= "000000";
				when "000101010000111110" => data <= "000000";
				when "000101010000111111" => data <= "000000";
				when "000101010001000000" => data <= "000000";
				when "000101010001000001" => data <= "000000";
				when "000101010001000010" => data <= "000000";
				when "000101010001000011" => data <= "000000";
				when "000101010001000100" => data <= "000000";
				when "000101010001000101" => data <= "000000";
				when "000101010001000110" => data <= "000000";
				when "000101010001000111" => data <= "000000";
				when "000101010001001000" => data <= "000000";
				when "000101010001001001" => data <= "000000";
				when "000101010001001010" => data <= "000000";
				when "000101010001001011" => data <= "000000";
				when "000101010001001100" => data <= "000000";
				when "000101010001001101" => data <= "000000";
				when "000101010001001110" => data <= "000000";
				when "000101010001001111" => data <= "000000";
				when "000101010001010000" => data <= "000000";
				when "000101010001010001" => data <= "000000";
				when "000101010001010010" => data <= "000000";
				when "000101010001010011" => data <= "000000";
				when "000101010001010100" => data <= "000000";
				when "000101010001010101" => data <= "000000";
				when "000101010001010110" => data <= "000000";
				when "000101010001010111" => data <= "000000";
				when "000101010001011000" => data <= "000000";
				when "000101010001011001" => data <= "000000";
				when "000101010001011010" => data <= "000000";
				when "000101010001011011" => data <= "000000";
				when "000101010001011100" => data <= "000000";
				when "000101010001011101" => data <= "000000";
				when "000101010001011110" => data <= "000000";
				when "000101010001011111" => data <= "000000";
				when "000101010001100000" => data <= "000000";
				when "000101010001100001" => data <= "000000";
				when "000101010001100010" => data <= "000000";
				when "000101010001100011" => data <= "000000";
				when "000101010001100100" => data <= "000000";
				when "000101010001100101" => data <= "000000";
				when "000101010001100110" => data <= "000000";
				when "000101010001100111" => data <= "000000";
				when "000101010001101000" => data <= "000000";
				when "000101010001101001" => data <= "000000";
				when "000101010001101010" => data <= "000000";
				when "000101010001101011" => data <= "000000";
				when "000101010001101100" => data <= "000000";
				when "000101010001101101" => data <= "000000";
				when "000101010001101110" => data <= "000000";
				when "000101010001101111" => data <= "000000";
				when "000101010001110000" => data <= "000000";
				when "000101010001110001" => data <= "000000";
				when "000101010001110010" => data <= "000000";
				when "000101010001110011" => data <= "000000";
				when "000101010001110100" => data <= "000000";
				when "000101010001110101" => data <= "000000";
				when "000101010001110110" => data <= "000000";
				when "000101010001110111" => data <= "000000";
				when "000101010001111000" => data <= "000000";
				when "000101010001111001" => data <= "000000";
				when "000101010001111010" => data <= "000000";
				when "000101010001111011" => data <= "000000";
				when "000101010001111100" => data <= "000000";
				when "000101010001111101" => data <= "000000";
				when "000101010001111110" => data <= "000000";
				when "000101010001111111" => data <= "000000";
				when "000101010010000000" => data <= "000000";
				when "000101010010000001" => data <= "000000";
				when "000101010010000010" => data <= "000000";
				when "000101010010000011" => data <= "000000";
				when "000101010010000100" => data <= "000000";
				when "000101010010000101" => data <= "000000";
				when "000101010010000110" => data <= "000000";
				when "000101010010000111" => data <= "000000";
				when "000101010010001000" => data <= "000000";
				when "000101010010001001" => data <= "000000";
				when "000101010010001010" => data <= "000000";
				when "000101010010001011" => data <= "000000";
				when "000101010010001100" => data <= "000000";
				when "000101010010001101" => data <= "000000";
				when "000101010010001110" => data <= "000000";
				when "000101010010001111" => data <= "000000";
				when "000101010010010000" => data <= "000000";
				when "000101010010010001" => data <= "000000";
				when "000101010010010010" => data <= "000000";
				when "000101010010010011" => data <= "000000";
				when "000101010010010100" => data <= "000000";
				when "000101010010010101" => data <= "000000";
				when "000101010010010110" => data <= "000000";
				when "000101010010010111" => data <= "000000";
				when "000101010010011000" => data <= "000000";
				when "000101010010011001" => data <= "000000";
				when "000101010010011010" => data <= "000000";
				when "000101010010011011" => data <= "000000";
				when "000101010010011100" => data <= "000000";
				when "000101010010011101" => data <= "000000";
				when "000101010010011110" => data <= "000000";
				when "000101010010011111" => data <= "000000";
				when "000101011000000000" => data <= "000000";
				when "000101011000000001" => data <= "000000";
				when "000101011000000010" => data <= "000000";
				when "000101011000000011" => data <= "000000";
				when "000101011000000100" => data <= "000000";
				when "000101011000000101" => data <= "000000";
				when "000101011000000110" => data <= "000000";
				when "000101011000000111" => data <= "000000";
				when "000101011000001000" => data <= "000000";
				when "000101011000001001" => data <= "000000";
				when "000101011000001010" => data <= "000000";
				when "000101011000001011" => data <= "000000";
				when "000101011000001100" => data <= "000000";
				when "000101011000001101" => data <= "000000";
				when "000101011000001110" => data <= "000000";
				when "000101011000001111" => data <= "000000";
				when "000101011000010000" => data <= "000000";
				when "000101011000010001" => data <= "000000";
				when "000101011000010010" => data <= "000000";
				when "000101011000010011" => data <= "000000";
				when "000101011000010100" => data <= "000000";
				when "000101011000010101" => data <= "000000";
				when "000101011000010110" => data <= "000000";
				when "000101011000010111" => data <= "000000";
				when "000101011000011000" => data <= "000000";
				when "000101011000011001" => data <= "000000";
				when "000101011000011010" => data <= "000000";
				when "000101011000011011" => data <= "000000";
				when "000101011000011100" => data <= "000000";
				when "000101011000011101" => data <= "000000";
				when "000101011000011110" => data <= "000000";
				when "000101011000011111" => data <= "000000";
				when "000101011000100000" => data <= "000000";
				when "000101011000100001" => data <= "000000";
				when "000101011000100010" => data <= "000000";
				when "000101011000100011" => data <= "000000";
				when "000101011000100100" => data <= "000000";
				when "000101011000100101" => data <= "000000";
				when "000101011000100110" => data <= "000000";
				when "000101011000100111" => data <= "000000";
				when "000101011000101000" => data <= "000000";
				when "000101011000101001" => data <= "000000";
				when "000101011000101010" => data <= "000000";
				when "000101011000101011" => data <= "000000";
				when "000101011000101100" => data <= "000000";
				when "000101011000101101" => data <= "000000";
				when "000101011000101110" => data <= "000000";
				when "000101011000101111" => data <= "000000";
				when "000101011000110000" => data <= "000000";
				when "000101011000110001" => data <= "000000";
				when "000101011000110010" => data <= "000000";
				when "000101011000110011" => data <= "000000";
				when "000101011000110100" => data <= "000000";
				when "000101011000110101" => data <= "000000";
				when "000101011000110110" => data <= "000000";
				when "000101011000110111" => data <= "000000";
				when "000101011000111000" => data <= "000000";
				when "000101011000111001" => data <= "000000";
				when "000101011000111010" => data <= "000000";
				when "000101011000111011" => data <= "000000";
				when "000101011000111100" => data <= "000000";
				when "000101011000111101" => data <= "000000";
				when "000101011000111110" => data <= "000000";
				when "000101011000111111" => data <= "000000";
				when "000101011001000000" => data <= "000000";
				when "000101011001000001" => data <= "000000";
				when "000101011001000010" => data <= "000000";
				when "000101011001000011" => data <= "000000";
				when "000101011001000100" => data <= "000000";
				when "000101011001000101" => data <= "000000";
				when "000101011001000110" => data <= "000000";
				when "000101011001000111" => data <= "000000";
				when "000101011001001000" => data <= "000000";
				when "000101011001001001" => data <= "000000";
				when "000101011001001010" => data <= "000000";
				when "000101011001001011" => data <= "000000";
				when "000101011001001100" => data <= "000000";
				when "000101011001001101" => data <= "000000";
				when "000101011001001110" => data <= "000000";
				when "000101011001001111" => data <= "000000";
				when "000101011001010000" => data <= "000000";
				when "000101011001010001" => data <= "000000";
				when "000101011001010010" => data <= "000000";
				when "000101011001010011" => data <= "000000";
				when "000101011001010100" => data <= "000000";
				when "000101011001010101" => data <= "000000";
				when "000101011001010110" => data <= "000000";
				when "000101011001010111" => data <= "000000";
				when "000101011001011000" => data <= "000000";
				when "000101011001011001" => data <= "000000";
				when "000101011001011010" => data <= "000000";
				when "000101011001011011" => data <= "000000";
				when "000101011001011100" => data <= "000000";
				when "000101011001011101" => data <= "000000";
				when "000101011001011110" => data <= "000000";
				when "000101011001011111" => data <= "000000";
				when "000101011001100000" => data <= "000000";
				when "000101011001100001" => data <= "000000";
				when "000101011001100010" => data <= "000000";
				when "000101011001100011" => data <= "000000";
				when "000101011001100100" => data <= "000000";
				when "000101011001100101" => data <= "000000";
				when "000101011001100110" => data <= "000000";
				when "000101011001100111" => data <= "000000";
				when "000101011001101000" => data <= "000000";
				when "000101011001101001" => data <= "000000";
				when "000101011001101010" => data <= "000000";
				when "000101011001101011" => data <= "000000";
				when "000101011001101100" => data <= "000000";
				when "000101011001101101" => data <= "000000";
				when "000101011001101110" => data <= "000000";
				when "000101011001101111" => data <= "000000";
				when "000101011001110000" => data <= "000000";
				when "000101011001110001" => data <= "000000";
				when "000101011001110010" => data <= "000000";
				when "000101011001110011" => data <= "000000";
				when "000101011001110100" => data <= "000000";
				when "000101011001110101" => data <= "000000";
				when "000101011001110110" => data <= "000000";
				when "000101011001110111" => data <= "000000";
				when "000101011001111000" => data <= "000000";
				when "000101011001111001" => data <= "000000";
				when "000101011001111010" => data <= "000000";
				when "000101011001111011" => data <= "000000";
				when "000101011001111100" => data <= "000000";
				when "000101011001111101" => data <= "000000";
				when "000101011001111110" => data <= "000000";
				when "000101011001111111" => data <= "000000";
				when "000101011010000000" => data <= "000000";
				when "000101011010000001" => data <= "000000";
				when "000101011010000010" => data <= "000000";
				when "000101011010000011" => data <= "000000";
				when "000101011010000100" => data <= "000000";
				when "000101011010000101" => data <= "000000";
				when "000101011010000110" => data <= "000000";
				when "000101011010000111" => data <= "000000";
				when "000101011010001000" => data <= "000000";
				when "000101011010001001" => data <= "000000";
				when "000101011010001010" => data <= "000000";
				when "000101011010001011" => data <= "000000";
				when "000101011010001100" => data <= "000000";
				when "000101011010001101" => data <= "000000";
				when "000101011010001110" => data <= "000000";
				when "000101011010001111" => data <= "000000";
				when "000101011010010000" => data <= "000000";
				when "000101011010010001" => data <= "000000";
				when "000101011010010010" => data <= "000000";
				when "000101011010010011" => data <= "000000";
				when "000101011010010100" => data <= "000000";
				when "000101011010010101" => data <= "000000";
				when "000101011010010110" => data <= "000000";
				when "000101011010010111" => data <= "000000";
				when "000101011010011000" => data <= "000000";
				when "000101011010011001" => data <= "000000";
				when "000101011010011010" => data <= "000000";
				when "000101011010011011" => data <= "000000";
				when "000101011010011100" => data <= "000000";
				when "000101011010011101" => data <= "000000";
				when "000101011010011110" => data <= "000000";
				when "000101011010011111" => data <= "000000";
				when "000101100000000000" => data <= "000000";
				when "000101100000000001" => data <= "000000";
				when "000101100000000010" => data <= "000000";
				when "000101100000000011" => data <= "000000";
				when "000101100000000100" => data <= "000000";
				when "000101100000000101" => data <= "000000";
				when "000101100000000110" => data <= "000000";
				when "000101100000000111" => data <= "000000";
				when "000101100000001000" => data <= "000000";
				when "000101100000001001" => data <= "000000";
				when "000101100000001010" => data <= "000000";
				when "000101100000001011" => data <= "000000";
				when "000101100000001100" => data <= "000000";
				when "000101100000001101" => data <= "000000";
				when "000101100000001110" => data <= "000000";
				when "000101100000001111" => data <= "000000";
				when "000101100000010000" => data <= "000000";
				when "000101100000010001" => data <= "000000";
				when "000101100000010010" => data <= "000000";
				when "000101100000010011" => data <= "000000";
				when "000101100000010100" => data <= "000000";
				when "000101100000010101" => data <= "000000";
				when "000101100000010110" => data <= "000000";
				when "000101100000010111" => data <= "000000";
				when "000101100000011000" => data <= "000000";
				when "000101100000011001" => data <= "000000";
				when "000101100000011010" => data <= "000000";
				when "000101100000011011" => data <= "000000";
				when "000101100000011100" => data <= "000000";
				when "000101100000011101" => data <= "000000";
				when "000101100000011110" => data <= "000000";
				when "000101100000011111" => data <= "000000";
				when "000101100000100000" => data <= "000000";
				when "000101100000100001" => data <= "000000";
				when "000101100000100010" => data <= "000000";
				when "000101100000100011" => data <= "000000";
				when "000101100000100100" => data <= "000000";
				when "000101100000100101" => data <= "000000";
				when "000101100000100110" => data <= "000000";
				when "000101100000100111" => data <= "000000";
				when "000101100000101000" => data <= "000000";
				when "000101100000101001" => data <= "000000";
				when "000101100000101010" => data <= "000000";
				when "000101100000101011" => data <= "000000";
				when "000101100000101100" => data <= "000000";
				when "000101100000101101" => data <= "000000";
				when "000101100000101110" => data <= "000000";
				when "000101100000101111" => data <= "000000";
				when "000101100000110000" => data <= "000000";
				when "000101100000110001" => data <= "000000";
				when "000101100000110010" => data <= "000000";
				when "000101100000110011" => data <= "000000";
				when "000101100000110100" => data <= "000000";
				when "000101100000110101" => data <= "000000";
				when "000101100000110110" => data <= "000000";
				when "000101100000110111" => data <= "000000";
				when "000101100000111000" => data <= "000000";
				when "000101100000111001" => data <= "000000";
				when "000101100000111010" => data <= "000000";
				when "000101100000111011" => data <= "000000";
				when "000101100000111100" => data <= "000000";
				when "000101100000111101" => data <= "000000";
				when "000101100000111110" => data <= "000000";
				when "000101100000111111" => data <= "000000";
				when "000101100001000000" => data <= "000000";
				when "000101100001000001" => data <= "000000";
				when "000101100001000010" => data <= "000000";
				when "000101100001000011" => data <= "000000";
				when "000101100001000100" => data <= "000000";
				when "000101100001000101" => data <= "000000";
				when "000101100001000110" => data <= "000000";
				when "000101100001000111" => data <= "000000";
				when "000101100001001000" => data <= "000000";
				when "000101100001001001" => data <= "000000";
				when "000101100001001010" => data <= "000000";
				when "000101100001001011" => data <= "000000";
				when "000101100001001100" => data <= "000000";
				when "000101100001001101" => data <= "000000";
				when "000101100001001110" => data <= "000000";
				when "000101100001001111" => data <= "000000";
				when "000101100001010000" => data <= "000000";
				when "000101100001010001" => data <= "000000";
				when "000101100001010010" => data <= "000000";
				when "000101100001010011" => data <= "000000";
				when "000101100001010100" => data <= "000000";
				when "000101100001010101" => data <= "000000";
				when "000101100001010110" => data <= "000000";
				when "000101100001010111" => data <= "000000";
				when "000101100001011000" => data <= "000000";
				when "000101100001011001" => data <= "000000";
				when "000101100001011010" => data <= "000000";
				when "000101100001011011" => data <= "000000";
				when "000101100001011100" => data <= "000000";
				when "000101100001011101" => data <= "000000";
				when "000101100001011110" => data <= "000000";
				when "000101100001011111" => data <= "000000";
				when "000101100001100000" => data <= "000000";
				when "000101100001100001" => data <= "000000";
				when "000101100001100010" => data <= "000000";
				when "000101100001100011" => data <= "000000";
				when "000101100001100100" => data <= "000000";
				when "000101100001100101" => data <= "000000";
				when "000101100001100110" => data <= "000000";
				when "000101100001100111" => data <= "000000";
				when "000101100001101000" => data <= "000000";
				when "000101100001101001" => data <= "000000";
				when "000101100001101010" => data <= "000000";
				when "000101100001101011" => data <= "000000";
				when "000101100001101100" => data <= "000000";
				when "000101100001101101" => data <= "000000";
				when "000101100001101110" => data <= "000000";
				when "000101100001101111" => data <= "000000";
				when "000101100001110000" => data <= "000000";
				when "000101100001110001" => data <= "000000";
				when "000101100001110010" => data <= "000000";
				when "000101100001110011" => data <= "000000";
				when "000101100001110100" => data <= "000000";
				when "000101100001110101" => data <= "000000";
				when "000101100001110110" => data <= "000000";
				when "000101100001110111" => data <= "000000";
				when "000101100001111000" => data <= "000000";
				when "000101100001111001" => data <= "000000";
				when "000101100001111010" => data <= "000000";
				when "000101100001111011" => data <= "000000";
				when "000101100001111100" => data <= "000000";
				when "000101100001111101" => data <= "000000";
				when "000101100001111110" => data <= "000000";
				when "000101100001111111" => data <= "000000";
				when "000101100010000000" => data <= "000000";
				when "000101100010000001" => data <= "000000";
				when "000101100010000010" => data <= "000000";
				when "000101100010000011" => data <= "000000";
				when "000101100010000100" => data <= "000000";
				when "000101100010000101" => data <= "000000";
				when "000101100010000110" => data <= "000000";
				when "000101100010000111" => data <= "000000";
				when "000101100010001000" => data <= "000000";
				when "000101100010001001" => data <= "000000";
				when "000101100010001010" => data <= "000000";
				when "000101100010001011" => data <= "000000";
				when "000101100010001100" => data <= "000000";
				when "000101100010001101" => data <= "000000";
				when "000101100010001110" => data <= "000000";
				when "000101100010001111" => data <= "000000";
				when "000101100010010000" => data <= "000000";
				when "000101100010010001" => data <= "000000";
				when "000101100010010010" => data <= "000000";
				when "000101100010010011" => data <= "000000";
				when "000101100010010100" => data <= "000000";
				when "000101100010010101" => data <= "000000";
				when "000101100010010110" => data <= "000000";
				when "000101100010010111" => data <= "000000";
				when "000101100010011000" => data <= "000000";
				when "000101100010011001" => data <= "000000";
				when "000101100010011010" => data <= "000000";
				when "000101100010011011" => data <= "000000";
				when "000101100010011100" => data <= "000000";
				when "000101100010011101" => data <= "000000";
				when "000101100010011110" => data <= "000000";
				when "000101100010011111" => data <= "000000";
				when "000101101000000000" => data <= "000000";
				when "000101101000000001" => data <= "000000";
				when "000101101000000010" => data <= "000000";
				when "000101101000000011" => data <= "000000";
				when "000101101000000100" => data <= "000000";
				when "000101101000000101" => data <= "000000";
				when "000101101000000110" => data <= "000000";
				when "000101101000000111" => data <= "000000";
				when "000101101000001000" => data <= "000000";
				when "000101101000001001" => data <= "000000";
				when "000101101000001010" => data <= "000000";
				when "000101101000001011" => data <= "000000";
				when "000101101000001100" => data <= "000000";
				when "000101101000001101" => data <= "000000";
				when "000101101000001110" => data <= "000000";
				when "000101101000001111" => data <= "000000";
				when "000101101000010000" => data <= "000000";
				when "000101101000010001" => data <= "000000";
				when "000101101000010010" => data <= "000000";
				when "000101101000010011" => data <= "000000";
				when "000101101000010100" => data <= "000000";
				when "000101101000010101" => data <= "000000";
				when "000101101000010110" => data <= "000000";
				when "000101101000010111" => data <= "000000";
				when "000101101000011000" => data <= "000000";
				when "000101101000011001" => data <= "000000";
				when "000101101000011010" => data <= "000000";
				when "000101101000011011" => data <= "000000";
				when "000101101000011100" => data <= "000000";
				when "000101101000011101" => data <= "000000";
				when "000101101000011110" => data <= "000000";
				when "000101101000011111" => data <= "000000";
				when "000101101000100000" => data <= "000000";
				when "000101101000100001" => data <= "000000";
				when "000101101000100010" => data <= "000000";
				when "000101101000100011" => data <= "000000";
				when "000101101000100100" => data <= "000000";
				when "000101101000100101" => data <= "000000";
				when "000101101000100110" => data <= "000000";
				when "000101101000100111" => data <= "000000";
				when "000101101000101000" => data <= "000000";
				when "000101101000101001" => data <= "000000";
				when "000101101000101010" => data <= "000000";
				when "000101101000101011" => data <= "000000";
				when "000101101000101100" => data <= "000000";
				when "000101101000101101" => data <= "000000";
				when "000101101000101110" => data <= "000000";
				when "000101101000101111" => data <= "000000";
				when "000101101000110000" => data <= "000000";
				when "000101101000110001" => data <= "000000";
				when "000101101000110010" => data <= "000000";
				when "000101101000110011" => data <= "000000";
				when "000101101000110100" => data <= "000000";
				when "000101101000110101" => data <= "000000";
				when "000101101000110110" => data <= "000000";
				when "000101101000110111" => data <= "000000";
				when "000101101000111000" => data <= "000000";
				when "000101101000111001" => data <= "000000";
				when "000101101000111010" => data <= "000000";
				when "000101101000111011" => data <= "000000";
				when "000101101000111100" => data <= "000000";
				when "000101101000111101" => data <= "000000";
				when "000101101000111110" => data <= "000000";
				when "000101101000111111" => data <= "000000";
				when "000101101001000000" => data <= "000000";
				when "000101101001000001" => data <= "000000";
				when "000101101001000010" => data <= "000000";
				when "000101101001000011" => data <= "000000";
				when "000101101001000100" => data <= "000000";
				when "000101101001000101" => data <= "000000";
				when "000101101001000110" => data <= "000000";
				when "000101101001000111" => data <= "000000";
				when "000101101001001000" => data <= "000000";
				when "000101101001001001" => data <= "000000";
				when "000101101001001010" => data <= "000000";
				when "000101101001001011" => data <= "000000";
				when "000101101001001100" => data <= "000000";
				when "000101101001001101" => data <= "000000";
				when "000101101001001110" => data <= "000000";
				when "000101101001001111" => data <= "000000";
				when "000101101001010000" => data <= "000000";
				when "000101101001010001" => data <= "000000";
				when "000101101001010010" => data <= "000000";
				when "000101101001010011" => data <= "000000";
				when "000101101001010100" => data <= "000000";
				when "000101101001010101" => data <= "000000";
				when "000101101001010110" => data <= "000000";
				when "000101101001010111" => data <= "000000";
				when "000101101001011000" => data <= "000000";
				when "000101101001011001" => data <= "000000";
				when "000101101001011010" => data <= "000000";
				when "000101101001011011" => data <= "000000";
				when "000101101001011100" => data <= "000000";
				when "000101101001011101" => data <= "000000";
				when "000101101001011110" => data <= "000000";
				when "000101101001011111" => data <= "000000";
				when "000101101001100000" => data <= "000000";
				when "000101101001100001" => data <= "000000";
				when "000101101001100010" => data <= "000000";
				when "000101101001100011" => data <= "000000";
				when "000101101001100100" => data <= "000000";
				when "000101101001100101" => data <= "000000";
				when "000101101001100110" => data <= "000000";
				when "000101101001100111" => data <= "000000";
				when "000101101001101000" => data <= "000000";
				when "000101101001101001" => data <= "000000";
				when "000101101001101010" => data <= "000000";
				when "000101101001101011" => data <= "000000";
				when "000101101001101100" => data <= "000000";
				when "000101101001101101" => data <= "000000";
				when "000101101001101110" => data <= "000000";
				when "000101101001101111" => data <= "000000";
				when "000101101001110000" => data <= "000000";
				when "000101101001110001" => data <= "000000";
				when "000101101001110010" => data <= "000000";
				when "000101101001110011" => data <= "000000";
				when "000101101001110100" => data <= "000000";
				when "000101101001110101" => data <= "000000";
				when "000101101001110110" => data <= "000000";
				when "000101101001110111" => data <= "000000";
				when "000101101001111000" => data <= "000000";
				when "000101101001111001" => data <= "000000";
				when "000101101001111010" => data <= "000000";
				when "000101101001111011" => data <= "000000";
				when "000101101001111100" => data <= "000000";
				when "000101101001111101" => data <= "000000";
				when "000101101001111110" => data <= "000000";
				when "000101101001111111" => data <= "000000";
				when "000101101010000000" => data <= "000000";
				when "000101101010000001" => data <= "000000";
				when "000101101010000010" => data <= "000000";
				when "000101101010000011" => data <= "000000";
				when "000101101010000100" => data <= "000000";
				when "000101101010000101" => data <= "000000";
				when "000101101010000110" => data <= "000000";
				when "000101101010000111" => data <= "000000";
				when "000101101010001000" => data <= "000000";
				when "000101101010001001" => data <= "000000";
				when "000101101010001010" => data <= "000000";
				when "000101101010001011" => data <= "000000";
				when "000101101010001100" => data <= "000000";
				when "000101101010001101" => data <= "000000";
				when "000101101010001110" => data <= "000000";
				when "000101101010001111" => data <= "000000";
				when "000101101010010000" => data <= "000000";
				when "000101101010010001" => data <= "000000";
				when "000101101010010010" => data <= "000000";
				when "000101101010010011" => data <= "000000";
				when "000101101010010100" => data <= "000000";
				when "000101101010010101" => data <= "000000";
				when "000101101010010110" => data <= "000000";
				when "000101101010010111" => data <= "000000";
				when "000101101010011000" => data <= "000000";
				when "000101101010011001" => data <= "000000";
				when "000101101010011010" => data <= "000000";
				when "000101101010011011" => data <= "000000";
				when "000101101010011100" => data <= "000000";
				when "000101101010011101" => data <= "000000";
				when "000101101010011110" => data <= "000000";
				when "000101101010011111" => data <= "000000";
				when "000101110000000000" => data <= "000000";
				when "000101110000000001" => data <= "000000";
				when "000101110000000010" => data <= "000000";
				when "000101110000000011" => data <= "000000";
				when "000101110000000100" => data <= "000000";
				when "000101110000000101" => data <= "000000";
				when "000101110000000110" => data <= "000000";
				when "000101110000000111" => data <= "000000";
				when "000101110000001000" => data <= "000000";
				when "000101110000001001" => data <= "000000";
				when "000101110000001010" => data <= "000000";
				when "000101110000001011" => data <= "000000";
				when "000101110000001100" => data <= "000000";
				when "000101110000001101" => data <= "000000";
				when "000101110000001110" => data <= "000000";
				when "000101110000001111" => data <= "000000";
				when "000101110000010000" => data <= "000000";
				when "000101110000010001" => data <= "000000";
				when "000101110000010010" => data <= "000000";
				when "000101110000010011" => data <= "000000";
				when "000101110000010100" => data <= "000000";
				when "000101110000010101" => data <= "000000";
				when "000101110000010110" => data <= "000000";
				when "000101110000010111" => data <= "000000";
				when "000101110000011000" => data <= "000000";
				when "000101110000011001" => data <= "000000";
				when "000101110000011010" => data <= "000000";
				when "000101110000011011" => data <= "000000";
				when "000101110000011100" => data <= "000000";
				when "000101110000011101" => data <= "000000";
				when "000101110000011110" => data <= "000000";
				when "000101110000011111" => data <= "000000";
				when "000101110000100000" => data <= "000000";
				when "000101110000100001" => data <= "000000";
				when "000101110000100010" => data <= "000000";
				when "000101110000100011" => data <= "000000";
				when "000101110000100100" => data <= "000000";
				when "000101110000100101" => data <= "000000";
				when "000101110000100110" => data <= "000000";
				when "000101110000100111" => data <= "000000";
				when "000101110000101000" => data <= "000000";
				when "000101110000101001" => data <= "000000";
				when "000101110000101010" => data <= "000000";
				when "000101110000101011" => data <= "000000";
				when "000101110000101100" => data <= "000000";
				when "000101110000101101" => data <= "000000";
				when "000101110000101110" => data <= "000000";
				when "000101110000101111" => data <= "000000";
				when "000101110000110000" => data <= "000000";
				when "000101110000110001" => data <= "000000";
				when "000101110000110010" => data <= "000000";
				when "000101110000110011" => data <= "000000";
				when "000101110000110100" => data <= "000000";
				when "000101110000110101" => data <= "000000";
				when "000101110000110110" => data <= "000000";
				when "000101110000110111" => data <= "000000";
				when "000101110000111000" => data <= "000000";
				when "000101110000111001" => data <= "000000";
				when "000101110000111010" => data <= "000000";
				when "000101110000111011" => data <= "000000";
				when "000101110000111100" => data <= "000000";
				when "000101110000111101" => data <= "000000";
				when "000101110000111110" => data <= "000000";
				when "000101110000111111" => data <= "000000";
				when "000101110001000000" => data <= "000000";
				when "000101110001000001" => data <= "000000";
				when "000101110001000010" => data <= "000000";
				when "000101110001000011" => data <= "000000";
				when "000101110001000100" => data <= "000000";
				when "000101110001000101" => data <= "000000";
				when "000101110001000110" => data <= "000000";
				when "000101110001000111" => data <= "000000";
				when "000101110001001000" => data <= "000000";
				when "000101110001001001" => data <= "000000";
				when "000101110001001010" => data <= "000000";
				when "000101110001001011" => data <= "000000";
				when "000101110001001100" => data <= "000000";
				when "000101110001001101" => data <= "000000";
				when "000101110001001110" => data <= "000000";
				when "000101110001001111" => data <= "000000";
				when "000101110001010000" => data <= "000000";
				when "000101110001010001" => data <= "000000";
				when "000101110001010010" => data <= "000000";
				when "000101110001010011" => data <= "000000";
				when "000101110001010100" => data <= "000000";
				when "000101110001010101" => data <= "000000";
				when "000101110001010110" => data <= "000000";
				when "000101110001010111" => data <= "000000";
				when "000101110001011000" => data <= "000000";
				when "000101110001011001" => data <= "000000";
				when "000101110001011010" => data <= "000000";
				when "000101110001011011" => data <= "000000";
				when "000101110001011100" => data <= "000000";
				when "000101110001011101" => data <= "000000";
				when "000101110001011110" => data <= "000000";
				when "000101110001011111" => data <= "000000";
				when "000101110001100000" => data <= "000000";
				when "000101110001100001" => data <= "000000";
				when "000101110001100010" => data <= "000000";
				when "000101110001100011" => data <= "000000";
				when "000101110001100100" => data <= "000000";
				when "000101110001100101" => data <= "000000";
				when "000101110001100110" => data <= "000000";
				when "000101110001100111" => data <= "000000";
				when "000101110001101000" => data <= "000000";
				when "000101110001101001" => data <= "000000";
				when "000101110001101010" => data <= "000000";
				when "000101110001101011" => data <= "000000";
				when "000101110001101100" => data <= "000000";
				when "000101110001101101" => data <= "000000";
				when "000101110001101110" => data <= "000000";
				when "000101110001101111" => data <= "000000";
				when "000101110001110000" => data <= "000000";
				when "000101110001110001" => data <= "000000";
				when "000101110001110010" => data <= "000000";
				when "000101110001110011" => data <= "000000";
				when "000101110001110100" => data <= "000000";
				when "000101110001110101" => data <= "000000";
				when "000101110001110110" => data <= "000000";
				when "000101110001110111" => data <= "000000";
				when "000101110001111000" => data <= "000000";
				when "000101110001111001" => data <= "000000";
				when "000101110001111010" => data <= "000000";
				when "000101110001111011" => data <= "000000";
				when "000101110001111100" => data <= "000000";
				when "000101110001111101" => data <= "000000";
				when "000101110001111110" => data <= "000000";
				when "000101110001111111" => data <= "000000";
				when "000101110010000000" => data <= "000000";
				when "000101110010000001" => data <= "000000";
				when "000101110010000010" => data <= "000000";
				when "000101110010000011" => data <= "000000";
				when "000101110010000100" => data <= "000000";
				when "000101110010000101" => data <= "000000";
				when "000101110010000110" => data <= "000000";
				when "000101110010000111" => data <= "000000";
				when "000101110010001000" => data <= "000000";
				when "000101110010001001" => data <= "000000";
				when "000101110010001010" => data <= "000000";
				when "000101110010001011" => data <= "000000";
				when "000101110010001100" => data <= "000000";
				when "000101110010001101" => data <= "000000";
				when "000101110010001110" => data <= "000000";
				when "000101110010001111" => data <= "000000";
				when "000101110010010000" => data <= "000000";
				when "000101110010010001" => data <= "000000";
				when "000101110010010010" => data <= "000000";
				when "000101110010010011" => data <= "000000";
				when "000101110010010100" => data <= "000000";
				when "000101110010010101" => data <= "000000";
				when "000101110010010110" => data <= "000000";
				when "000101110010010111" => data <= "000000";
				when "000101110010011000" => data <= "000000";
				when "000101110010011001" => data <= "000000";
				when "000101110010011010" => data <= "000000";
				when "000101110010011011" => data <= "000000";
				when "000101110010011100" => data <= "000000";
				when "000101110010011101" => data <= "000000";
				when "000101110010011110" => data <= "000000";
				when "000101110010011111" => data <= "000000";
				when "000101111000000000" => data <= "000000";
				when "000101111000000001" => data <= "000000";
				when "000101111000000010" => data <= "000000";
				when "000101111000000011" => data <= "000000";
				when "000101111000000100" => data <= "000000";
				when "000101111000000101" => data <= "000000";
				when "000101111000000110" => data <= "000000";
				when "000101111000000111" => data <= "000000";
				when "000101111000001000" => data <= "000000";
				when "000101111000001001" => data <= "000000";
				when "000101111000001010" => data <= "000000";
				when "000101111000001011" => data <= "000000";
				when "000101111000001100" => data <= "000000";
				when "000101111000001101" => data <= "000000";
				when "000101111000001110" => data <= "000000";
				when "000101111000001111" => data <= "000000";
				when "000101111000010000" => data <= "000000";
				when "000101111000010001" => data <= "000000";
				when "000101111000010010" => data <= "000000";
				when "000101111000010011" => data <= "000000";
				when "000101111000010100" => data <= "000000";
				when "000101111000010101" => data <= "000000";
				when "000101111000010110" => data <= "000000";
				when "000101111000010111" => data <= "000000";
				when "000101111000011000" => data <= "000000";
				when "000101111000011001" => data <= "000000";
				when "000101111000011010" => data <= "000000";
				when "000101111000011011" => data <= "000000";
				when "000101111000011100" => data <= "000000";
				when "000101111000011101" => data <= "000000";
				when "000101111000011110" => data <= "000000";
				when "000101111000011111" => data <= "000000";
				when "000101111000100000" => data <= "000000";
				when "000101111000100001" => data <= "000000";
				when "000101111000100010" => data <= "000000";
				when "000101111000100011" => data <= "000000";
				when "000101111000100100" => data <= "000000";
				when "000101111000100101" => data <= "000000";
				when "000101111000100110" => data <= "000000";
				when "000101111000100111" => data <= "000000";
				when "000101111000101000" => data <= "000000";
				when "000101111000101001" => data <= "000000";
				when "000101111000101010" => data <= "000000";
				when "000101111000101011" => data <= "000000";
				when "000101111000101100" => data <= "000000";
				when "000101111000101101" => data <= "000000";
				when "000101111000101110" => data <= "000000";
				when "000101111000101111" => data <= "000000";
				when "000101111000110000" => data <= "000000";
				when "000101111000110001" => data <= "000000";
				when "000101111000110010" => data <= "000000";
				when "000101111000110011" => data <= "000000";
				when "000101111000110100" => data <= "000000";
				when "000101111000110101" => data <= "000000";
				when "000101111000110110" => data <= "000000";
				when "000101111000110111" => data <= "000000";
				when "000101111000111000" => data <= "000000";
				when "000101111000111001" => data <= "000000";
				when "000101111000111010" => data <= "000000";
				when "000101111000111011" => data <= "000000";
				when "000101111000111100" => data <= "000000";
				when "000101111000111101" => data <= "000000";
				when "000101111000111110" => data <= "000000";
				when "000101111000111111" => data <= "000000";
				when "000101111001000000" => data <= "000000";
				when "000101111001000001" => data <= "000000";
				when "000101111001000010" => data <= "000000";
				when "000101111001000011" => data <= "000000";
				when "000101111001000100" => data <= "000000";
				when "000101111001000101" => data <= "000000";
				when "000101111001000110" => data <= "000000";
				when "000101111001000111" => data <= "000000";
				when "000101111001001000" => data <= "000000";
				when "000101111001001001" => data <= "000000";
				when "000101111001001010" => data <= "000000";
				when "000101111001001011" => data <= "000000";
				when "000101111001001100" => data <= "000000";
				when "000101111001001101" => data <= "000000";
				when "000101111001001110" => data <= "000000";
				when "000101111001001111" => data <= "000000";
				when "000101111001010000" => data <= "000000";
				when "000101111001010001" => data <= "000000";
				when "000101111001010010" => data <= "000000";
				when "000101111001010011" => data <= "000000";
				when "000101111001010100" => data <= "000000";
				when "000101111001010101" => data <= "000000";
				when "000101111001010110" => data <= "000000";
				when "000101111001010111" => data <= "000000";
				when "000101111001011000" => data <= "000000";
				when "000101111001011001" => data <= "000000";
				when "000101111001011010" => data <= "000000";
				when "000101111001011011" => data <= "000000";
				when "000101111001011100" => data <= "000000";
				when "000101111001011101" => data <= "000000";
				when "000101111001011110" => data <= "000000";
				when "000101111001011111" => data <= "000000";
				when "000101111001100000" => data <= "000000";
				when "000101111001100001" => data <= "000000";
				when "000101111001100010" => data <= "000000";
				when "000101111001100011" => data <= "000000";
				when "000101111001100100" => data <= "000000";
				when "000101111001100101" => data <= "000000";
				when "000101111001100110" => data <= "000000";
				when "000101111001100111" => data <= "000000";
				when "000101111001101000" => data <= "000000";
				when "000101111001101001" => data <= "000000";
				when "000101111001101010" => data <= "000000";
				when "000101111001101011" => data <= "000000";
				when "000101111001101100" => data <= "000000";
				when "000101111001101101" => data <= "000000";
				when "000101111001101110" => data <= "000000";
				when "000101111001101111" => data <= "000000";
				when "000101111001110000" => data <= "000000";
				when "000101111001110001" => data <= "000000";
				when "000101111001110010" => data <= "000000";
				when "000101111001110011" => data <= "000000";
				when "000101111001110100" => data <= "000000";
				when "000101111001110101" => data <= "000000";
				when "000101111001110110" => data <= "000000";
				when "000101111001110111" => data <= "000000";
				when "000101111001111000" => data <= "000000";
				when "000101111001111001" => data <= "000000";
				when "000101111001111010" => data <= "000000";
				when "000101111001111011" => data <= "000000";
				when "000101111001111100" => data <= "000000";
				when "000101111001111101" => data <= "000000";
				when "000101111001111110" => data <= "000000";
				when "000101111001111111" => data <= "000000";
				when "000101111010000000" => data <= "000000";
				when "000101111010000001" => data <= "000000";
				when "000101111010000010" => data <= "000000";
				when "000101111010000011" => data <= "000000";
				when "000101111010000100" => data <= "000000";
				when "000101111010000101" => data <= "000000";
				when "000101111010000110" => data <= "000000";
				when "000101111010000111" => data <= "000000";
				when "000101111010001000" => data <= "000000";
				when "000101111010001001" => data <= "000000";
				when "000101111010001010" => data <= "000000";
				when "000101111010001011" => data <= "000000";
				when "000101111010001100" => data <= "000000";
				when "000101111010001101" => data <= "000000";
				when "000101111010001110" => data <= "000000";
				when "000101111010001111" => data <= "000000";
				when "000101111010010000" => data <= "000000";
				when "000101111010010001" => data <= "000000";
				when "000101111010010010" => data <= "000000";
				when "000101111010010011" => data <= "000000";
				when "000101111010010100" => data <= "000000";
				when "000101111010010101" => data <= "000000";
				when "000101111010010110" => data <= "000000";
				when "000101111010010111" => data <= "000000";
				when "000101111010011000" => data <= "000000";
				when "000101111010011001" => data <= "000000";
				when "000101111010011010" => data <= "000000";
				when "000101111010011011" => data <= "000000";
				when "000101111010011100" => data <= "000000";
				when "000101111010011101" => data <= "000000";
				when "000101111010011110" => data <= "000000";
				when "000101111010011111" => data <= "000000";
				when "000110000000000000" => data <= "000000";
				when "000110000000000001" => data <= "000000";
				when "000110000000000010" => data <= "000000";
				when "000110000000000011" => data <= "000000";
				when "000110000000000100" => data <= "000000";
				when "000110000000000101" => data <= "000000";
				when "000110000000000110" => data <= "000000";
				when "000110000000000111" => data <= "000000";
				when "000110000000001000" => data <= "000000";
				when "000110000000001001" => data <= "000000";
				when "000110000000001010" => data <= "000000";
				when "000110000000001011" => data <= "000000";
				when "000110000000001100" => data <= "000000";
				when "000110000000001101" => data <= "000000";
				when "000110000000001110" => data <= "000000";
				when "000110000000001111" => data <= "000000";
				when "000110000000010000" => data <= "000000";
				when "000110000000010001" => data <= "000000";
				when "000110000000010010" => data <= "000000";
				when "000110000000010011" => data <= "000000";
				when "000110000000010100" => data <= "000000";
				when "000110000000010101" => data <= "000000";
				when "000110000000010110" => data <= "000000";
				when "000110000000010111" => data <= "000000";
				when "000110000000011000" => data <= "000000";
				when "000110000000011001" => data <= "000000";
				when "000110000000011010" => data <= "000000";
				when "000110000000011011" => data <= "000000";
				when "000110000000011100" => data <= "000000";
				when "000110000000011101" => data <= "000000";
				when "000110000000011110" => data <= "000000";
				when "000110000000011111" => data <= "000000";
				when "000110000000100000" => data <= "000000";
				when "000110000000100001" => data <= "000000";
				when "000110000000100010" => data <= "000000";
				when "000110000000100011" => data <= "000000";
				when "000110000000100100" => data <= "000000";
				when "000110000000100101" => data <= "000000";
				when "000110000000100110" => data <= "000000";
				when "000110000000100111" => data <= "000000";
				when "000110000000101000" => data <= "000000";
				when "000110000000101001" => data <= "000000";
				when "000110000000101010" => data <= "000000";
				when "000110000000101011" => data <= "000000";
				when "000110000000101100" => data <= "000000";
				when "000110000000101101" => data <= "000000";
				when "000110000000101110" => data <= "000000";
				when "000110000000101111" => data <= "000000";
				when "000110000000110000" => data <= "000000";
				when "000110000000110001" => data <= "000000";
				when "000110000000110010" => data <= "000000";
				when "000110000000110011" => data <= "000000";
				when "000110000000110100" => data <= "000000";
				when "000110000000110101" => data <= "000000";
				when "000110000000110110" => data <= "000000";
				when "000110000000110111" => data <= "000000";
				when "000110000000111000" => data <= "000000";
				when "000110000000111001" => data <= "000000";
				when "000110000000111010" => data <= "000000";
				when "000110000000111011" => data <= "000000";
				when "000110000000111100" => data <= "000000";
				when "000110000000111101" => data <= "000000";
				when "000110000000111110" => data <= "000000";
				when "000110000000111111" => data <= "000000";
				when "000110000001000000" => data <= "000000";
				when "000110000001000001" => data <= "000000";
				when "000110000001000010" => data <= "000000";
				when "000110000001000011" => data <= "000000";
				when "000110000001000100" => data <= "000000";
				when "000110000001000101" => data <= "000000";
				when "000110000001000110" => data <= "000000";
				when "000110000001000111" => data <= "000000";
				when "000110000001001000" => data <= "000000";
				when "000110000001001001" => data <= "000000";
				when "000110000001001010" => data <= "000000";
				when "000110000001001011" => data <= "000000";
				when "000110000001001100" => data <= "000000";
				when "000110000001001101" => data <= "000000";
				when "000110000001001110" => data <= "000000";
				when "000110000001001111" => data <= "000000";
				when "000110000001010000" => data <= "000000";
				when "000110000001010001" => data <= "000000";
				when "000110000001010010" => data <= "000000";
				when "000110000001010011" => data <= "000000";
				when "000110000001010100" => data <= "000000";
				when "000110000001010101" => data <= "000000";
				when "000110000001010110" => data <= "000000";
				when "000110000001010111" => data <= "000000";
				when "000110000001011000" => data <= "000000";
				when "000110000001011001" => data <= "000000";
				when "000110000001011010" => data <= "000000";
				when "000110000001011011" => data <= "000000";
				when "000110000001011100" => data <= "000000";
				when "000110000001011101" => data <= "000000";
				when "000110000001011110" => data <= "000000";
				when "000110000001011111" => data <= "000000";
				when "000110000001100000" => data <= "000000";
				when "000110000001100001" => data <= "000000";
				when "000110000001100010" => data <= "000000";
				when "000110000001100011" => data <= "000000";
				when "000110000001100100" => data <= "000000";
				when "000110000001100101" => data <= "000000";
				when "000110000001100110" => data <= "000000";
				when "000110000001100111" => data <= "000000";
				when "000110000001101000" => data <= "000000";
				when "000110000001101001" => data <= "000000";
				when "000110000001101010" => data <= "000000";
				when "000110000001101011" => data <= "000000";
				when "000110000001101100" => data <= "000000";
				when "000110000001101101" => data <= "000000";
				when "000110000001101110" => data <= "000000";
				when "000110000001101111" => data <= "000000";
				when "000110000001110000" => data <= "000000";
				when "000110000001110001" => data <= "000000";
				when "000110000001110010" => data <= "000000";
				when "000110000001110011" => data <= "000000";
				when "000110000001110100" => data <= "000000";
				when "000110000001110101" => data <= "000000";
				when "000110000001110110" => data <= "000000";
				when "000110000001110111" => data <= "000000";
				when "000110000001111000" => data <= "000000";
				when "000110000001111001" => data <= "000000";
				when "000110000001111010" => data <= "000000";
				when "000110000001111011" => data <= "000000";
				when "000110000001111100" => data <= "000000";
				when "000110000001111101" => data <= "000000";
				when "000110000001111110" => data <= "000000";
				when "000110000001111111" => data <= "000000";
				when "000110000010000000" => data <= "000000";
				when "000110000010000001" => data <= "000000";
				when "000110000010000010" => data <= "000000";
				when "000110000010000011" => data <= "000000";
				when "000110000010000100" => data <= "000000";
				when "000110000010000101" => data <= "000000";
				when "000110000010000110" => data <= "000000";
				when "000110000010000111" => data <= "000000";
				when "000110000010001000" => data <= "000000";
				when "000110000010001001" => data <= "000000";
				when "000110000010001010" => data <= "000000";
				when "000110000010001011" => data <= "000000";
				when "000110000010001100" => data <= "000000";
				when "000110000010001101" => data <= "000000";
				when "000110000010001110" => data <= "000000";
				when "000110000010001111" => data <= "000000";
				when "000110000010010000" => data <= "000000";
				when "000110000010010001" => data <= "000000";
				when "000110000010010010" => data <= "000000";
				when "000110000010010011" => data <= "000000";
				when "000110000010010100" => data <= "000000";
				when "000110000010010101" => data <= "000000";
				when "000110000010010110" => data <= "000000";
				when "000110000010010111" => data <= "000000";
				when "000110000010011000" => data <= "000000";
				when "000110000010011001" => data <= "000000";
				when "000110000010011010" => data <= "000000";
				when "000110000010011011" => data <= "000000";
				when "000110000010011100" => data <= "000000";
				when "000110000010011101" => data <= "000000";
				when "000110000010011110" => data <= "000000";
				when "000110000010011111" => data <= "000000";
				when "000110001000000000" => data <= "000000";
				when "000110001000000001" => data <= "000000";
				when "000110001000000010" => data <= "000000";
				when "000110001000000011" => data <= "000000";
				when "000110001000000100" => data <= "000000";
				when "000110001000000101" => data <= "000000";
				when "000110001000000110" => data <= "000000";
				when "000110001000000111" => data <= "000000";
				when "000110001000001000" => data <= "000000";
				when "000110001000001001" => data <= "000000";
				when "000110001000001010" => data <= "000000";
				when "000110001000001011" => data <= "000000";
				when "000110001000001100" => data <= "000000";
				when "000110001000001101" => data <= "000000";
				when "000110001000001110" => data <= "000000";
				when "000110001000001111" => data <= "000000";
				when "000110001000010000" => data <= "000000";
				when "000110001000010001" => data <= "000000";
				when "000110001000010010" => data <= "000000";
				when "000110001000010011" => data <= "000000";
				when "000110001000010100" => data <= "000000";
				when "000110001000010101" => data <= "000000";
				when "000110001000010110" => data <= "000000";
				when "000110001000010111" => data <= "000000";
				when "000110001000011000" => data <= "000000";
				when "000110001000011001" => data <= "000000";
				when "000110001000011010" => data <= "000000";
				when "000110001000011011" => data <= "000000";
				when "000110001000011100" => data <= "000000";
				when "000110001000011101" => data <= "000000";
				when "000110001000011110" => data <= "000000";
				when "000110001000011111" => data <= "000000";
				when "000110001000100000" => data <= "000000";
				when "000110001000100001" => data <= "000000";
				when "000110001000100010" => data <= "000000";
				when "000110001000100011" => data <= "000000";
				when "000110001000100100" => data <= "000000";
				when "000110001000100101" => data <= "000000";
				when "000110001000100110" => data <= "000000";
				when "000110001000100111" => data <= "000000";
				when "000110001000101000" => data <= "000000";
				when "000110001000101001" => data <= "000000";
				when "000110001000101010" => data <= "000000";
				when "000110001000101011" => data <= "000000";
				when "000110001000101100" => data <= "000000";
				when "000110001000101101" => data <= "000000";
				when "000110001000101110" => data <= "000000";
				when "000110001000101111" => data <= "000000";
				when "000110001000110000" => data <= "000000";
				when "000110001000110001" => data <= "000000";
				when "000110001000110010" => data <= "000000";
				when "000110001000110011" => data <= "000000";
				when "000110001000110100" => data <= "000000";
				when "000110001000110101" => data <= "000000";
				when "000110001000110110" => data <= "000000";
				when "000110001000110111" => data <= "000000";
				when "000110001000111000" => data <= "000000";
				when "000110001000111001" => data <= "000000";
				when "000110001000111010" => data <= "000000";
				when "000110001000111011" => data <= "000000";
				when "000110001000111100" => data <= "000000";
				when "000110001000111101" => data <= "000000";
				when "000110001000111110" => data <= "000000";
				when "000110001000111111" => data <= "000000";
				when "000110001001000000" => data <= "000000";
				when "000110001001000001" => data <= "000000";
				when "000110001001000010" => data <= "000000";
				when "000110001001000011" => data <= "000000";
				when "000110001001000100" => data <= "000000";
				when "000110001001000101" => data <= "000000";
				when "000110001001000110" => data <= "000000";
				when "000110001001000111" => data <= "000000";
				when "000110001001001000" => data <= "000000";
				when "000110001001001001" => data <= "000000";
				when "000110001001001010" => data <= "000000";
				when "000110001001001011" => data <= "000000";
				when "000110001001001100" => data <= "000000";
				when "000110001001001101" => data <= "000000";
				when "000110001001001110" => data <= "000000";
				when "000110001001001111" => data <= "000000";
				when "000110001001010000" => data <= "000000";
				when "000110001001010001" => data <= "000000";
				when "000110001001010010" => data <= "000000";
				when "000110001001010011" => data <= "000000";
				when "000110001001010100" => data <= "000000";
				when "000110001001010101" => data <= "000000";
				when "000110001001010110" => data <= "000000";
				when "000110001001010111" => data <= "000000";
				when "000110001001011000" => data <= "000000";
				when "000110001001011001" => data <= "000000";
				when "000110001001011010" => data <= "000000";
				when "000110001001011011" => data <= "000000";
				when "000110001001011100" => data <= "000000";
				when "000110001001011101" => data <= "000000";
				when "000110001001011110" => data <= "000000";
				when "000110001001011111" => data <= "000000";
				when "000110001001100000" => data <= "000000";
				when "000110001001100001" => data <= "000000";
				when "000110001001100010" => data <= "000000";
				when "000110001001100011" => data <= "000000";
				when "000110001001100100" => data <= "000000";
				when "000110001001100101" => data <= "000000";
				when "000110001001100110" => data <= "000000";
				when "000110001001100111" => data <= "000000";
				when "000110001001101000" => data <= "000000";
				when "000110001001101001" => data <= "000000";
				when "000110001001101010" => data <= "000000";
				when "000110001001101011" => data <= "000000";
				when "000110001001101100" => data <= "000000";
				when "000110001001101101" => data <= "000000";
				when "000110001001101110" => data <= "000000";
				when "000110001001101111" => data <= "000000";
				when "000110001001110000" => data <= "000000";
				when "000110001001110001" => data <= "000000";
				when "000110001001110010" => data <= "000000";
				when "000110001001110011" => data <= "000000";
				when "000110001001110100" => data <= "000000";
				when "000110001001110101" => data <= "000000";
				when "000110001001110110" => data <= "000000";
				when "000110001001110111" => data <= "000000";
				when "000110001001111000" => data <= "000000";
				when "000110001001111001" => data <= "000000";
				when "000110001001111010" => data <= "000000";
				when "000110001001111011" => data <= "000000";
				when "000110001001111100" => data <= "000000";
				when "000110001001111101" => data <= "000000";
				when "000110001001111110" => data <= "000000";
				when "000110001001111111" => data <= "000000";
				when "000110001010000000" => data <= "000000";
				when "000110001010000001" => data <= "000000";
				when "000110001010000010" => data <= "000000";
				when "000110001010000011" => data <= "000000";
				when "000110001010000100" => data <= "000000";
				when "000110001010000101" => data <= "000000";
				when "000110001010000110" => data <= "000000";
				when "000110001010000111" => data <= "000000";
				when "000110001010001000" => data <= "000000";
				when "000110001010001001" => data <= "000000";
				when "000110001010001010" => data <= "000000";
				when "000110001010001011" => data <= "000000";
				when "000110001010001100" => data <= "000000";
				when "000110001010001101" => data <= "000000";
				when "000110001010001110" => data <= "000000";
				when "000110001010001111" => data <= "000000";
				when "000110001010010000" => data <= "000000";
				when "000110001010010001" => data <= "000000";
				when "000110001010010010" => data <= "000000";
				when "000110001010010011" => data <= "000000";
				when "000110001010010100" => data <= "000000";
				when "000110001010010101" => data <= "000000";
				when "000110001010010110" => data <= "000000";
				when "000110001010010111" => data <= "000000";
				when "000110001010011000" => data <= "000000";
				when "000110001010011001" => data <= "000000";
				when "000110001010011010" => data <= "000000";
				when "000110001010011011" => data <= "000000";
				when "000110001010011100" => data <= "000000";
				when "000110001010011101" => data <= "000000";
				when "000110001010011110" => data <= "000000";
				when "000110001010011111" => data <= "000000";
				when "000110010000000000" => data <= "000000";
				when "000110010000000001" => data <= "000000";
				when "000110010000000010" => data <= "000000";
				when "000110010000000011" => data <= "000000";
				when "000110010000000100" => data <= "000000";
				when "000110010000000101" => data <= "000000";
				when "000110010000000110" => data <= "000000";
				when "000110010000000111" => data <= "000000";
				when "000110010000001000" => data <= "000000";
				when "000110010000001001" => data <= "000000";
				when "000110010000001010" => data <= "000000";
				when "000110010000001011" => data <= "000000";
				when "000110010000001100" => data <= "000000";
				when "000110010000001101" => data <= "000000";
				when "000110010000001110" => data <= "000000";
				when "000110010000001111" => data <= "000000";
				when "000110010000010000" => data <= "000000";
				when "000110010000010001" => data <= "000000";
				when "000110010000010010" => data <= "000000";
				when "000110010000010011" => data <= "000000";
				when "000110010000010100" => data <= "000000";
				when "000110010000010101" => data <= "000000";
				when "000110010000010110" => data <= "000000";
				when "000110010000010111" => data <= "000000";
				when "000110010000011000" => data <= "000000";
				when "000110010000011001" => data <= "000000";
				when "000110010000011010" => data <= "000000";
				when "000110010000011011" => data <= "000000";
				when "000110010000011100" => data <= "000000";
				when "000110010000011101" => data <= "000000";
				when "000110010000011110" => data <= "000000";
				when "000110010000011111" => data <= "000000";
				when "000110010000100000" => data <= "000000";
				when "000110010000100001" => data <= "000000";
				when "000110010000100010" => data <= "000000";
				when "000110010000100011" => data <= "000000";
				when "000110010000100100" => data <= "000000";
				when "000110010000100101" => data <= "000000";
				when "000110010000100110" => data <= "000000";
				when "000110010000100111" => data <= "000000";
				when "000110010000101000" => data <= "000000";
				when "000110010000101001" => data <= "000000";
				when "000110010000101010" => data <= "000000";
				when "000110010000101011" => data <= "000000";
				when "000110010000101100" => data <= "000000";
				when "000110010000101101" => data <= "000000";
				when "000110010000101110" => data <= "000000";
				when "000110010000101111" => data <= "000000";
				when "000110010000110000" => data <= "000000";
				when "000110010000110001" => data <= "000000";
				when "000110010000110010" => data <= "000000";
				when "000110010000110011" => data <= "000000";
				when "000110010000110100" => data <= "000000";
				when "000110010000110101" => data <= "000000";
				when "000110010000110110" => data <= "000000";
				when "000110010000110111" => data <= "000000";
				when "000110010000111000" => data <= "000000";
				when "000110010000111001" => data <= "000000";
				when "000110010000111010" => data <= "000000";
				when "000110010000111011" => data <= "000000";
				when "000110010000111100" => data <= "000000";
				when "000110010000111101" => data <= "000000";
				when "000110010000111110" => data <= "000000";
				when "000110010000111111" => data <= "000000";
				when "000110010001000000" => data <= "000000";
				when "000110010001000001" => data <= "000000";
				when "000110010001000010" => data <= "000000";
				when "000110010001000011" => data <= "000000";
				when "000110010001000100" => data <= "000000";
				when "000110010001000101" => data <= "000000";
				when "000110010001000110" => data <= "000000";
				when "000110010001000111" => data <= "000000";
				when "000110010001001000" => data <= "000000";
				when "000110010001001001" => data <= "000000";
				when "000110010001001010" => data <= "000000";
				when "000110010001001011" => data <= "000000";
				when "000110010001001100" => data <= "000000";
				when "000110010001001101" => data <= "000000";
				when "000110010001001110" => data <= "000000";
				when "000110010001001111" => data <= "000000";
				when "000110010001010000" => data <= "000000";
				when "000110010001010001" => data <= "000000";
				when "000110010001010010" => data <= "000000";
				when "000110010001010011" => data <= "000000";
				when "000110010001010100" => data <= "000000";
				when "000110010001010101" => data <= "000000";
				when "000110010001010110" => data <= "000000";
				when "000110010001010111" => data <= "000000";
				when "000110010001011000" => data <= "000000";
				when "000110010001011001" => data <= "000000";
				when "000110010001011010" => data <= "000000";
				when "000110010001011011" => data <= "000000";
				when "000110010001011100" => data <= "000000";
				when "000110010001011101" => data <= "000000";
				when "000110010001011110" => data <= "000000";
				when "000110010001011111" => data <= "000000";
				when "000110010001100000" => data <= "000000";
				when "000110010001100001" => data <= "000000";
				when "000110010001100010" => data <= "000000";
				when "000110010001100011" => data <= "000000";
				when "000110010001100100" => data <= "000000";
				when "000110010001100101" => data <= "000000";
				when "000110010001100110" => data <= "000000";
				when "000110010001100111" => data <= "000000";
				when "000110010001101000" => data <= "000000";
				when "000110010001101001" => data <= "000000";
				when "000110010001101010" => data <= "000000";
				when "000110010001101011" => data <= "000000";
				when "000110010001101100" => data <= "000000";
				when "000110010001101101" => data <= "000000";
				when "000110010001101110" => data <= "000000";
				when "000110010001101111" => data <= "000000";
				when "000110010001110000" => data <= "000000";
				when "000110010001110001" => data <= "000000";
				when "000110010001110010" => data <= "000000";
				when "000110010001110011" => data <= "000000";
				when "000110010001110100" => data <= "000000";
				when "000110010001110101" => data <= "000000";
				when "000110010001110110" => data <= "000000";
				when "000110010001110111" => data <= "000000";
				when "000110010001111000" => data <= "000000";
				when "000110010001111001" => data <= "000000";
				when "000110010001111010" => data <= "000000";
				when "000110010001111011" => data <= "000000";
				when "000110010001111100" => data <= "000000";
				when "000110010001111101" => data <= "000000";
				when "000110010001111110" => data <= "000000";
				when "000110010001111111" => data <= "000000";
				when "000110010010000000" => data <= "000000";
				when "000110010010000001" => data <= "000000";
				when "000110010010000010" => data <= "000000";
				when "000110010010000011" => data <= "000000";
				when "000110010010000100" => data <= "000000";
				when "000110010010000101" => data <= "000000";
				when "000110010010000110" => data <= "000000";
				when "000110010010000111" => data <= "000000";
				when "000110010010001000" => data <= "000000";
				when "000110010010001001" => data <= "000000";
				when "000110010010001010" => data <= "000000";
				when "000110010010001011" => data <= "000000";
				when "000110010010001100" => data <= "000000";
				when "000110010010001101" => data <= "000000";
				when "000110010010001110" => data <= "000000";
				when "000110010010001111" => data <= "000000";
				when "000110010010010000" => data <= "000000";
				when "000110010010010001" => data <= "000000";
				when "000110010010010010" => data <= "000000";
				when "000110010010010011" => data <= "000000";
				when "000110010010010100" => data <= "000000";
				when "000110010010010101" => data <= "000000";
				when "000110010010010110" => data <= "000000";
				when "000110010010010111" => data <= "000000";
				when "000110010010011000" => data <= "000000";
				when "000110010010011001" => data <= "000000";
				when "000110010010011010" => data <= "000000";
				when "000110010010011011" => data <= "000000";
				when "000110010010011100" => data <= "000000";
				when "000110010010011101" => data <= "000000";
				when "000110010010011110" => data <= "000000";
				when "000110010010011111" => data <= "000000";
				when "000110011000000000" => data <= "000000";
				when "000110011000000001" => data <= "000000";
				when "000110011000000010" => data <= "000000";
				when "000110011000000011" => data <= "000000";
				when "000110011000000100" => data <= "000000";
				when "000110011000000101" => data <= "000000";
				when "000110011000000110" => data <= "000000";
				when "000110011000000111" => data <= "000000";
				when "000110011000001000" => data <= "000000";
				when "000110011000001001" => data <= "000000";
				when "000110011000001010" => data <= "000000";
				when "000110011000001011" => data <= "000000";
				when "000110011000001100" => data <= "000000";
				when "000110011000001101" => data <= "000000";
				when "000110011000001110" => data <= "000000";
				when "000110011000001111" => data <= "000000";
				when "000110011000010000" => data <= "000000";
				when "000110011000010001" => data <= "000000";
				when "000110011000010010" => data <= "000000";
				when "000110011000010011" => data <= "000000";
				when "000110011000010100" => data <= "000000";
				when "000110011000010101" => data <= "000000";
				when "000110011000010110" => data <= "000000";
				when "000110011000010111" => data <= "000000";
				when "000110011000011000" => data <= "000000";
				when "000110011000011001" => data <= "000000";
				when "000110011000011010" => data <= "000000";
				when "000110011000011011" => data <= "000000";
				when "000110011000011100" => data <= "000000";
				when "000110011000011101" => data <= "000000";
				when "000110011000011110" => data <= "000000";
				when "000110011000011111" => data <= "000000";
				when "000110011000100000" => data <= "000000";
				when "000110011000100001" => data <= "000000";
				when "000110011000100010" => data <= "000000";
				when "000110011000100011" => data <= "000000";
				when "000110011000100100" => data <= "000000";
				when "000110011000100101" => data <= "000000";
				when "000110011000100110" => data <= "000000";
				when "000110011000100111" => data <= "000000";
				when "000110011000101000" => data <= "000000";
				when "000110011000101001" => data <= "000000";
				when "000110011000101010" => data <= "000000";
				when "000110011000101011" => data <= "000000";
				when "000110011000101100" => data <= "000000";
				when "000110011000101101" => data <= "000000";
				when "000110011000101110" => data <= "000000";
				when "000110011000101111" => data <= "000000";
				when "000110011000110000" => data <= "000000";
				when "000110011000110001" => data <= "000000";
				when "000110011000110010" => data <= "000000";
				when "000110011000110011" => data <= "000000";
				when "000110011000110100" => data <= "000000";
				when "000110011000110101" => data <= "000000";
				when "000110011000110110" => data <= "000000";
				when "000110011000110111" => data <= "000000";
				when "000110011000111000" => data <= "000000";
				when "000110011000111001" => data <= "000000";
				when "000110011000111010" => data <= "000000";
				when "000110011000111011" => data <= "000000";
				when "000110011000111100" => data <= "000000";
				when "000110011000111101" => data <= "000000";
				when "000110011000111110" => data <= "000000";
				when "000110011000111111" => data <= "000000";
				when "000110011001000000" => data <= "000000";
				when "000110011001000001" => data <= "000000";
				when "000110011001000010" => data <= "000000";
				when "000110011001000011" => data <= "000000";
				when "000110011001000100" => data <= "000000";
				when "000110011001000101" => data <= "000000";
				when "000110011001000110" => data <= "000000";
				when "000110011001000111" => data <= "000000";
				when "000110011001001000" => data <= "000000";
				when "000110011001001001" => data <= "000000";
				when "000110011001001010" => data <= "000000";
				when "000110011001001011" => data <= "000000";
				when "000110011001001100" => data <= "000000";
				when "000110011001001101" => data <= "000000";
				when "000110011001001110" => data <= "000000";
				when "000110011001001111" => data <= "000000";
				when "000110011001010000" => data <= "000000";
				when "000110011001010001" => data <= "000000";
				when "000110011001010010" => data <= "000000";
				when "000110011001010011" => data <= "000000";
				when "000110011001010100" => data <= "000000";
				when "000110011001010101" => data <= "000000";
				when "000110011001010110" => data <= "000000";
				when "000110011001010111" => data <= "000000";
				when "000110011001011000" => data <= "000000";
				when "000110011001011001" => data <= "000000";
				when "000110011001011010" => data <= "000000";
				when "000110011001011011" => data <= "000000";
				when "000110011001011100" => data <= "000000";
				when "000110011001011101" => data <= "000000";
				when "000110011001011110" => data <= "000000";
				when "000110011001011111" => data <= "000000";
				when "000110011001100000" => data <= "000000";
				when "000110011001100001" => data <= "000000";
				when "000110011001100010" => data <= "000000";
				when "000110011001100011" => data <= "000000";
				when "000110011001100100" => data <= "000000";
				when "000110011001100101" => data <= "000000";
				when "000110011001100110" => data <= "000000";
				when "000110011001100111" => data <= "000000";
				when "000110011001101000" => data <= "000000";
				when "000110011001101001" => data <= "000000";
				when "000110011001101010" => data <= "000000";
				when "000110011001101011" => data <= "000000";
				when "000110011001101100" => data <= "000000";
				when "000110011001101101" => data <= "000000";
				when "000110011001101110" => data <= "000000";
				when "000110011001101111" => data <= "000000";
				when "000110011001110000" => data <= "000000";
				when "000110011001110001" => data <= "000000";
				when "000110011001110010" => data <= "000000";
				when "000110011001110011" => data <= "000000";
				when "000110011001110100" => data <= "000000";
				when "000110011001110101" => data <= "000000";
				when "000110011001110110" => data <= "000000";
				when "000110011001110111" => data <= "000000";
				when "000110011001111000" => data <= "000000";
				when "000110011001111001" => data <= "000000";
				when "000110011001111010" => data <= "000000";
				when "000110011001111011" => data <= "000000";
				when "000110011001111100" => data <= "000000";
				when "000110011001111101" => data <= "000000";
				when "000110011001111110" => data <= "000000";
				when "000110011001111111" => data <= "000000";
				when "000110011010000000" => data <= "000000";
				when "000110011010000001" => data <= "000000";
				when "000110011010000010" => data <= "000000";
				when "000110011010000011" => data <= "000000";
				when "000110011010000100" => data <= "000000";
				when "000110011010000101" => data <= "000000";
				when "000110011010000110" => data <= "000000";
				when "000110011010000111" => data <= "000000";
				when "000110011010001000" => data <= "000000";
				when "000110011010001001" => data <= "000000";
				when "000110011010001010" => data <= "000000";
				when "000110011010001011" => data <= "000000";
				when "000110011010001100" => data <= "000000";
				when "000110011010001101" => data <= "000000";
				when "000110011010001110" => data <= "000000";
				when "000110011010001111" => data <= "000000";
				when "000110011010010000" => data <= "000000";
				when "000110011010010001" => data <= "000000";
				when "000110011010010010" => data <= "000000";
				when "000110011010010011" => data <= "000000";
				when "000110011010010100" => data <= "000000";
				when "000110011010010101" => data <= "000000";
				when "000110011010010110" => data <= "000000";
				when "000110011010010111" => data <= "000000";
				when "000110011010011000" => data <= "000000";
				when "000110011010011001" => data <= "000000";
				when "000110011010011010" => data <= "000000";
				when "000110011010011011" => data <= "000000";
				when "000110011010011100" => data <= "000000";
				when "000110011010011101" => data <= "000000";
				when "000110011010011110" => data <= "000000";
				when "000110011010011111" => data <= "000000";
				when "000110100000000000" => data <= "000000";
				when "000110100000000001" => data <= "000000";
				when "000110100000000010" => data <= "000000";
				when "000110100000000011" => data <= "000000";
				when "000110100000000100" => data <= "000000";
				when "000110100000000101" => data <= "000000";
				when "000110100000000110" => data <= "000000";
				when "000110100000000111" => data <= "000000";
				when "000110100000001000" => data <= "000000";
				when "000110100000001001" => data <= "000000";
				when "000110100000001010" => data <= "000000";
				when "000110100000001011" => data <= "000000";
				when "000110100000001100" => data <= "000000";
				when "000110100000001101" => data <= "000000";
				when "000110100000001110" => data <= "000000";
				when "000110100000001111" => data <= "000000";
				when "000110100000010000" => data <= "000000";
				when "000110100000010001" => data <= "000000";
				when "000110100000010010" => data <= "000000";
				when "000110100000010011" => data <= "000000";
				when "000110100000010100" => data <= "000000";
				when "000110100000010101" => data <= "000000";
				when "000110100000010110" => data <= "000000";
				when "000110100000010111" => data <= "000000";
				when "000110100000011000" => data <= "000000";
				when "000110100000011001" => data <= "000000";
				when "000110100000011010" => data <= "000000";
				when "000110100000011011" => data <= "000000";
				when "000110100000011100" => data <= "000000";
				when "000110100000011101" => data <= "000000";
				when "000110100000011110" => data <= "000000";
				when "000110100000011111" => data <= "000000";
				when "000110100000100000" => data <= "000000";
				when "000110100000100001" => data <= "000000";
				when "000110100000100010" => data <= "000000";
				when "000110100000100011" => data <= "000000";
				when "000110100000100100" => data <= "000000";
				when "000110100000100101" => data <= "000000";
				when "000110100000100110" => data <= "000000";
				when "000110100000100111" => data <= "000000";
				when "000110100000101000" => data <= "000000";
				when "000110100000101001" => data <= "000000";
				when "000110100000101010" => data <= "000000";
				when "000110100000101011" => data <= "000000";
				when "000110100000101100" => data <= "000000";
				when "000110100000101101" => data <= "000000";
				when "000110100000101110" => data <= "000000";
				when "000110100000101111" => data <= "000000";
				when "000110100000110000" => data <= "000000";
				when "000110100000110001" => data <= "000000";
				when "000110100000110010" => data <= "000000";
				when "000110100000110011" => data <= "000000";
				when "000110100000110100" => data <= "000000";
				when "000110100000110101" => data <= "000000";
				when "000110100000110110" => data <= "000000";
				when "000110100000110111" => data <= "000000";
				when "000110100000111000" => data <= "000000";
				when "000110100000111001" => data <= "000000";
				when "000110100000111010" => data <= "000000";
				when "000110100000111011" => data <= "000000";
				when "000110100000111100" => data <= "000000";
				when "000110100000111101" => data <= "000000";
				when "000110100000111110" => data <= "000000";
				when "000110100000111111" => data <= "000000";
				when "000110100001000000" => data <= "000000";
				when "000110100001000001" => data <= "000000";
				when "000110100001000010" => data <= "000000";
				when "000110100001000011" => data <= "000000";
				when "000110100001000100" => data <= "000000";
				when "000110100001000101" => data <= "000000";
				when "000110100001000110" => data <= "000000";
				when "000110100001000111" => data <= "000000";
				when "000110100001001000" => data <= "000000";
				when "000110100001001001" => data <= "000000";
				when "000110100001001010" => data <= "000000";
				when "000110100001001011" => data <= "000000";
				when "000110100001001100" => data <= "000000";
				when "000110100001001101" => data <= "000000";
				when "000110100001001110" => data <= "000000";
				when "000110100001001111" => data <= "000000";
				when "000110100001010000" => data <= "000000";
				when "000110100001010001" => data <= "000000";
				when "000110100001010010" => data <= "000000";
				when "000110100001010011" => data <= "000000";
				when "000110100001010100" => data <= "000000";
				when "000110100001010101" => data <= "000000";
				when "000110100001010110" => data <= "000000";
				when "000110100001010111" => data <= "000000";
				when "000110100001011000" => data <= "000000";
				when "000110100001011001" => data <= "000000";
				when "000110100001011010" => data <= "000000";
				when "000110100001011011" => data <= "000000";
				when "000110100001011100" => data <= "000000";
				when "000110100001011101" => data <= "000000";
				when "000110100001011110" => data <= "000000";
				when "000110100001011111" => data <= "000000";
				when "000110100001100000" => data <= "000000";
				when "000110100001100001" => data <= "000000";
				when "000110100001100010" => data <= "000000";
				when "000110100001100011" => data <= "000000";
				when "000110100001100100" => data <= "000000";
				when "000110100001100101" => data <= "000000";
				when "000110100001100110" => data <= "000000";
				when "000110100001100111" => data <= "000000";
				when "000110100001101000" => data <= "000000";
				when "000110100001101001" => data <= "000000";
				when "000110100001101010" => data <= "000000";
				when "000110100001101011" => data <= "000000";
				when "000110100001101100" => data <= "000000";
				when "000110100001101101" => data <= "000000";
				when "000110100001101110" => data <= "000000";
				when "000110100001101111" => data <= "000000";
				when "000110100001110000" => data <= "000000";
				when "000110100001110001" => data <= "000000";
				when "000110100001110010" => data <= "000000";
				when "000110100001110011" => data <= "000000";
				when "000110100001110100" => data <= "000000";
				when "000110100001110101" => data <= "000000";
				when "000110100001110110" => data <= "000000";
				when "000110100001110111" => data <= "000000";
				when "000110100001111000" => data <= "000000";
				when "000110100001111001" => data <= "000000";
				when "000110100001111010" => data <= "000000";
				when "000110100001111011" => data <= "000000";
				when "000110100001111100" => data <= "000000";
				when "000110100001111101" => data <= "000000";
				when "000110100001111110" => data <= "000000";
				when "000110100001111111" => data <= "000000";
				when "000110100010000000" => data <= "000000";
				when "000110100010000001" => data <= "000000";
				when "000110100010000010" => data <= "000000";
				when "000110100010000011" => data <= "000000";
				when "000110100010000100" => data <= "000000";
				when "000110100010000101" => data <= "000000";
				when "000110100010000110" => data <= "000000";
				when "000110100010000111" => data <= "000000";
				when "000110100010001000" => data <= "000000";
				when "000110100010001001" => data <= "000000";
				when "000110100010001010" => data <= "000000";
				when "000110100010001011" => data <= "000000";
				when "000110100010001100" => data <= "000000";
				when "000110100010001101" => data <= "000000";
				when "000110100010001110" => data <= "000000";
				when "000110100010001111" => data <= "000000";
				when "000110100010010000" => data <= "000000";
				when "000110100010010001" => data <= "000000";
				when "000110100010010010" => data <= "000000";
				when "000110100010010011" => data <= "000000";
				when "000110100010010100" => data <= "000000";
				when "000110100010010101" => data <= "000000";
				when "000110100010010110" => data <= "000000";
				when "000110100010010111" => data <= "000000";
				when "000110100010011000" => data <= "000000";
				when "000110100010011001" => data <= "000000";
				when "000110100010011010" => data <= "000000";
				when "000110100010011011" => data <= "000000";
				when "000110100010011100" => data <= "000000";
				when "000110100010011101" => data <= "000000";
				when "000110100010011110" => data <= "000000";
				when "000110100010011111" => data <= "000000";
				when "000110101000000000" => data <= "000000";
				when "000110101000000001" => data <= "000000";
				when "000110101000000010" => data <= "000000";
				when "000110101000000011" => data <= "000000";
				when "000110101000000100" => data <= "000000";
				when "000110101000000101" => data <= "000000";
				when "000110101000000110" => data <= "000000";
				when "000110101000000111" => data <= "000000";
				when "000110101000001000" => data <= "000000";
				when "000110101000001001" => data <= "000000";
				when "000110101000001010" => data <= "000000";
				when "000110101000001011" => data <= "000000";
				when "000110101000001100" => data <= "000000";
				when "000110101000001101" => data <= "000000";
				when "000110101000001110" => data <= "000000";
				when "000110101000001111" => data <= "000000";
				when "000110101000010000" => data <= "000000";
				when "000110101000010001" => data <= "000000";
				when "000110101000010010" => data <= "000000";
				when "000110101000010011" => data <= "000000";
				when "000110101000010100" => data <= "000000";
				when "000110101000010101" => data <= "000000";
				when "000110101000010110" => data <= "000000";
				when "000110101000010111" => data <= "000000";
				when "000110101000011000" => data <= "000000";
				when "000110101000011001" => data <= "000000";
				when "000110101000011010" => data <= "000000";
				when "000110101000011011" => data <= "000000";
				when "000110101000011100" => data <= "000000";
				when "000110101000011101" => data <= "000000";
				when "000110101000011110" => data <= "000000";
				when "000110101000011111" => data <= "000000";
				when "000110101000100000" => data <= "000000";
				when "000110101000100001" => data <= "000000";
				when "000110101000100010" => data <= "000000";
				when "000110101000100011" => data <= "000000";
				when "000110101000100100" => data <= "000000";
				when "000110101000100101" => data <= "000000";
				when "000110101000100110" => data <= "000000";
				when "000110101000100111" => data <= "000000";
				when "000110101000101000" => data <= "000000";
				when "000110101000101001" => data <= "000000";
				when "000110101000101010" => data <= "000000";
				when "000110101000101011" => data <= "000000";
				when "000110101000101100" => data <= "000000";
				when "000110101000101101" => data <= "000000";
				when "000110101000101110" => data <= "000000";
				when "000110101000101111" => data <= "000000";
				when "000110101000110000" => data <= "000000";
				when "000110101000110001" => data <= "000000";
				when "000110101000110010" => data <= "000000";
				when "000110101000110011" => data <= "000000";
				when "000110101000110100" => data <= "000000";
				when "000110101000110101" => data <= "000000";
				when "000110101000110110" => data <= "000000";
				when "000110101000110111" => data <= "000000";
				when "000110101000111000" => data <= "000000";
				when "000110101000111001" => data <= "000000";
				when "000110101000111010" => data <= "000000";
				when "000110101000111011" => data <= "000000";
				when "000110101000111100" => data <= "000000";
				when "000110101000111101" => data <= "000000";
				when "000110101000111110" => data <= "000000";
				when "000110101000111111" => data <= "000000";
				when "000110101001000000" => data <= "000000";
				when "000110101001000001" => data <= "000000";
				when "000110101001000010" => data <= "000000";
				when "000110101001000011" => data <= "000000";
				when "000110101001000100" => data <= "000000";
				when "000110101001000101" => data <= "000000";
				when "000110101001000110" => data <= "000000";
				when "000110101001000111" => data <= "000000";
				when "000110101001001000" => data <= "000000";
				when "000110101001001001" => data <= "000000";
				when "000110101001001010" => data <= "000000";
				when "000110101001001011" => data <= "000000";
				when "000110101001001100" => data <= "000000";
				when "000110101001001101" => data <= "000000";
				when "000110101001001110" => data <= "000000";
				when "000110101001001111" => data <= "000000";
				when "000110101001010000" => data <= "000000";
				when "000110101001010001" => data <= "000000";
				when "000110101001010010" => data <= "000000";
				when "000110101001010011" => data <= "000000";
				when "000110101001010100" => data <= "000000";
				when "000110101001010101" => data <= "000000";
				when "000110101001010110" => data <= "000000";
				when "000110101001010111" => data <= "000000";
				when "000110101001011000" => data <= "000000";
				when "000110101001011001" => data <= "000000";
				when "000110101001011010" => data <= "000000";
				when "000110101001011011" => data <= "000000";
				when "000110101001011100" => data <= "000000";
				when "000110101001011101" => data <= "000000";
				when "000110101001011110" => data <= "000000";
				when "000110101001011111" => data <= "000000";
				when "000110101001100000" => data <= "000000";
				when "000110101001100001" => data <= "000000";
				when "000110101001100010" => data <= "000000";
				when "000110101001100011" => data <= "000000";
				when "000110101001100100" => data <= "000000";
				when "000110101001100101" => data <= "000000";
				when "000110101001100110" => data <= "000000";
				when "000110101001100111" => data <= "000000";
				when "000110101001101000" => data <= "000000";
				when "000110101001101001" => data <= "000000";
				when "000110101001101010" => data <= "000000";
				when "000110101001101011" => data <= "000000";
				when "000110101001101100" => data <= "000000";
				when "000110101001101101" => data <= "000000";
				when "000110101001101110" => data <= "000000";
				when "000110101001101111" => data <= "000000";
				when "000110101001110000" => data <= "000000";
				when "000110101001110001" => data <= "000000";
				when "000110101001110010" => data <= "000000";
				when "000110101001110011" => data <= "000000";
				when "000110101001110100" => data <= "000000";
				when "000110101001110101" => data <= "000000";
				when "000110101001110110" => data <= "000000";
				when "000110101001110111" => data <= "000000";
				when "000110101001111000" => data <= "000000";
				when "000110101001111001" => data <= "000000";
				when "000110101001111010" => data <= "000000";
				when "000110101001111011" => data <= "000000";
				when "000110101001111100" => data <= "000000";
				when "000110101001111101" => data <= "000000";
				when "000110101001111110" => data <= "000000";
				when "000110101001111111" => data <= "000000";
				when "000110101010000000" => data <= "000000";
				when "000110101010000001" => data <= "000000";
				when "000110101010000010" => data <= "000000";
				when "000110101010000011" => data <= "000000";
				when "000110101010000100" => data <= "000000";
				when "000110101010000101" => data <= "000000";
				when "000110101010000110" => data <= "000000";
				when "000110101010000111" => data <= "000000";
				when "000110101010001000" => data <= "000000";
				when "000110101010001001" => data <= "000000";
				when "000110101010001010" => data <= "000000";
				when "000110101010001011" => data <= "000000";
				when "000110101010001100" => data <= "000000";
				when "000110101010001101" => data <= "000000";
				when "000110101010001110" => data <= "000000";
				when "000110101010001111" => data <= "000000";
				when "000110101010010000" => data <= "000000";
				when "000110101010010001" => data <= "000000";
				when "000110101010010010" => data <= "000000";
				when "000110101010010011" => data <= "000000";
				when "000110101010010100" => data <= "000000";
				when "000110101010010101" => data <= "000000";
				when "000110101010010110" => data <= "000000";
				when "000110101010010111" => data <= "000000";
				when "000110101010011000" => data <= "000000";
				when "000110101010011001" => data <= "000000";
				when "000110101010011010" => data <= "000000";
				when "000110101010011011" => data <= "000000";
				when "000110101010011100" => data <= "000000";
				when "000110101010011101" => data <= "000000";
				when "000110101010011110" => data <= "000000";
				when "000110101010011111" => data <= "000000";
				when "000110110000000000" => data <= "000000";
				when "000110110000000001" => data <= "000000";
				when "000110110000000010" => data <= "000000";
				when "000110110000000011" => data <= "000000";
				when "000110110000000100" => data <= "000000";
				when "000110110000000101" => data <= "000000";
				when "000110110000000110" => data <= "000000";
				when "000110110000000111" => data <= "000000";
				when "000110110000001000" => data <= "000000";
				when "000110110000001001" => data <= "000000";
				when "000110110000001010" => data <= "000000";
				when "000110110000001011" => data <= "000000";
				when "000110110000001100" => data <= "000000";
				when "000110110000001101" => data <= "000000";
				when "000110110000001110" => data <= "000000";
				when "000110110000001111" => data <= "000000";
				when "000110110000010000" => data <= "000000";
				when "000110110000010001" => data <= "000000";
				when "000110110000010010" => data <= "000000";
				when "000110110000010011" => data <= "000000";
				when "000110110000010100" => data <= "000000";
				when "000110110000010101" => data <= "000000";
				when "000110110000010110" => data <= "000000";
				when "000110110000010111" => data <= "000000";
				when "000110110000011000" => data <= "000000";
				when "000110110000011001" => data <= "000000";
				when "000110110000011010" => data <= "000000";
				when "000110110000011011" => data <= "000000";
				when "000110110000011100" => data <= "000000";
				when "000110110000011101" => data <= "000000";
				when "000110110000011110" => data <= "000000";
				when "000110110000011111" => data <= "000000";
				when "000110110000100000" => data <= "000000";
				when "000110110000100001" => data <= "000000";
				when "000110110000100010" => data <= "000000";
				when "000110110000100011" => data <= "000000";
				when "000110110000100100" => data <= "000000";
				when "000110110000100101" => data <= "000000";
				when "000110110000100110" => data <= "000000";
				when "000110110000100111" => data <= "000000";
				when "000110110000101000" => data <= "000000";
				when "000110110000101001" => data <= "000000";
				when "000110110000101010" => data <= "000000";
				when "000110110000101011" => data <= "000000";
				when "000110110000101100" => data <= "000000";
				when "000110110000101101" => data <= "000000";
				when "000110110000101110" => data <= "000000";
				when "000110110000101111" => data <= "000000";
				when "000110110000110000" => data <= "000000";
				when "000110110000110001" => data <= "000000";
				when "000110110000110010" => data <= "000000";
				when "000110110000110011" => data <= "000000";
				when "000110110000110100" => data <= "000000";
				when "000110110000110101" => data <= "000000";
				when "000110110000110110" => data <= "000000";
				when "000110110000110111" => data <= "000000";
				when "000110110000111000" => data <= "000000";
				when "000110110000111001" => data <= "000000";
				when "000110110000111010" => data <= "000000";
				when "000110110000111011" => data <= "000000";
				when "000110110000111100" => data <= "000000";
				when "000110110000111101" => data <= "000000";
				when "000110110000111110" => data <= "000000";
				when "000110110000111111" => data <= "000000";
				when "000110110001000000" => data <= "000000";
				when "000110110001000001" => data <= "000000";
				when "000110110001000010" => data <= "000000";
				when "000110110001000011" => data <= "000000";
				when "000110110001000100" => data <= "000000";
				when "000110110001000101" => data <= "000000";
				when "000110110001000110" => data <= "000000";
				when "000110110001000111" => data <= "000000";
				when "000110110001001000" => data <= "000000";
				when "000110110001001001" => data <= "000000";
				when "000110110001001010" => data <= "000000";
				when "000110110001001011" => data <= "000000";
				when "000110110001001100" => data <= "000000";
				when "000110110001001101" => data <= "000000";
				when "000110110001001110" => data <= "000000";
				when "000110110001001111" => data <= "000000";
				when "000110110001010000" => data <= "000000";
				when "000110110001010001" => data <= "000000";
				when "000110110001010010" => data <= "000000";
				when "000110110001010011" => data <= "000000";
				when "000110110001010100" => data <= "000000";
				when "000110110001010101" => data <= "000000";
				when "000110110001010110" => data <= "000000";
				when "000110110001010111" => data <= "000000";
				when "000110110001011000" => data <= "000000";
				when "000110110001011001" => data <= "000000";
				when "000110110001011010" => data <= "000000";
				when "000110110001011011" => data <= "000000";
				when "000110110001011100" => data <= "000000";
				when "000110110001011101" => data <= "000000";
				when "000110110001011110" => data <= "000000";
				when "000110110001011111" => data <= "000000";
				when "000110110001100000" => data <= "000000";
				when "000110110001100001" => data <= "000000";
				when "000110110001100010" => data <= "000000";
				when "000110110001100011" => data <= "000000";
				when "000110110001100100" => data <= "000000";
				when "000110110001100101" => data <= "000000";
				when "000110110001100110" => data <= "000000";
				when "000110110001100111" => data <= "000000";
				when "000110110001101000" => data <= "000000";
				when "000110110001101001" => data <= "000000";
				when "000110110001101010" => data <= "000000";
				when "000110110001101011" => data <= "000000";
				when "000110110001101100" => data <= "000000";
				when "000110110001101101" => data <= "000000";
				when "000110110001101110" => data <= "000000";
				when "000110110001101111" => data <= "000000";
				when "000110110001110000" => data <= "000000";
				when "000110110001110001" => data <= "000000";
				when "000110110001110010" => data <= "000000";
				when "000110110001110011" => data <= "000000";
				when "000110110001110100" => data <= "000000";
				when "000110110001110101" => data <= "000000";
				when "000110110001110110" => data <= "000000";
				when "000110110001110111" => data <= "000000";
				when "000110110001111000" => data <= "000000";
				when "000110110001111001" => data <= "000000";
				when "000110110001111010" => data <= "000000";
				when "000110110001111011" => data <= "000000";
				when "000110110001111100" => data <= "000000";
				when "000110110001111101" => data <= "000000";
				when "000110110001111110" => data <= "000000";
				when "000110110001111111" => data <= "000000";
				when "000110110010000000" => data <= "000000";
				when "000110110010000001" => data <= "000000";
				when "000110110010000010" => data <= "000000";
				when "000110110010000011" => data <= "000000";
				when "000110110010000100" => data <= "000000";
				when "000110110010000101" => data <= "000000";
				when "000110110010000110" => data <= "000000";
				when "000110110010000111" => data <= "000000";
				when "000110110010001000" => data <= "000000";
				when "000110110010001001" => data <= "000000";
				when "000110110010001010" => data <= "000000";
				when "000110110010001011" => data <= "000000";
				when "000110110010001100" => data <= "000000";
				when "000110110010001101" => data <= "000000";
				when "000110110010001110" => data <= "000000";
				when "000110110010001111" => data <= "000000";
				when "000110110010010000" => data <= "000000";
				when "000110110010010001" => data <= "000000";
				when "000110110010010010" => data <= "000000";
				when "000110110010010011" => data <= "000000";
				when "000110110010010100" => data <= "000000";
				when "000110110010010101" => data <= "000000";
				when "000110110010010110" => data <= "000000";
				when "000110110010010111" => data <= "000000";
				when "000110110010011000" => data <= "000000";
				when "000110110010011001" => data <= "000000";
				when "000110110010011010" => data <= "000000";
				when "000110110010011011" => data <= "000000";
				when "000110110010011100" => data <= "000000";
				when "000110110010011101" => data <= "000000";
				when "000110110010011110" => data <= "000000";
				when "000110110010011111" => data <= "000000";
				when "000110111000000000" => data <= "000000";
				when "000110111000000001" => data <= "000000";
				when "000110111000000010" => data <= "000000";
				when "000110111000000011" => data <= "000000";
				when "000110111000000100" => data <= "000000";
				when "000110111000000101" => data <= "000000";
				when "000110111000000110" => data <= "000000";
				when "000110111000000111" => data <= "000000";
				when "000110111000001000" => data <= "000000";
				when "000110111000001001" => data <= "000000";
				when "000110111000001010" => data <= "000000";
				when "000110111000001011" => data <= "000000";
				when "000110111000001100" => data <= "000000";
				when "000110111000001101" => data <= "000000";
				when "000110111000001110" => data <= "000000";
				when "000110111000001111" => data <= "000000";
				when "000110111000010000" => data <= "000000";
				when "000110111000010001" => data <= "000000";
				when "000110111000010010" => data <= "000000";
				when "000110111000010011" => data <= "000000";
				when "000110111000010100" => data <= "000000";
				when "000110111000010101" => data <= "000000";
				when "000110111000010110" => data <= "000000";
				when "000110111000010111" => data <= "000000";
				when "000110111000011000" => data <= "000000";
				when "000110111000011001" => data <= "000000";
				when "000110111000011010" => data <= "000000";
				when "000110111000011011" => data <= "000000";
				when "000110111000011100" => data <= "000000";
				when "000110111000011101" => data <= "000000";
				when "000110111000011110" => data <= "000000";
				when "000110111000011111" => data <= "000000";
				when "000110111000100000" => data <= "000000";
				when "000110111000100001" => data <= "000000";
				when "000110111000100010" => data <= "000000";
				when "000110111000100011" => data <= "000000";
				when "000110111000100100" => data <= "000000";
				when "000110111000100101" => data <= "000000";
				when "000110111000100110" => data <= "000000";
				when "000110111000100111" => data <= "000000";
				when "000110111000101000" => data <= "000000";
				when "000110111000101001" => data <= "000000";
				when "000110111000101010" => data <= "000000";
				when "000110111000101011" => data <= "000000";
				when "000110111000101100" => data <= "000000";
				when "000110111000101101" => data <= "000000";
				when "000110111000101110" => data <= "000000";
				when "000110111000101111" => data <= "000000";
				when "000110111000110000" => data <= "000000";
				when "000110111000110001" => data <= "000000";
				when "000110111000110010" => data <= "000000";
				when "000110111000110011" => data <= "000000";
				when "000110111000110100" => data <= "000000";
				when "000110111000110101" => data <= "000000";
				when "000110111000110110" => data <= "000000";
				when "000110111000110111" => data <= "000000";
				when "000110111000111000" => data <= "000000";
				when "000110111000111001" => data <= "000000";
				when "000110111000111010" => data <= "000000";
				when "000110111000111011" => data <= "000000";
				when "000110111000111100" => data <= "000000";
				when "000110111000111101" => data <= "000000";
				when "000110111000111110" => data <= "000000";
				when "000110111000111111" => data <= "000000";
				when "000110111001000000" => data <= "000000";
				when "000110111001000001" => data <= "000000";
				when "000110111001000010" => data <= "000000";
				when "000110111001000011" => data <= "000000";
				when "000110111001000100" => data <= "000000";
				when "000110111001000101" => data <= "000000";
				when "000110111001000110" => data <= "000000";
				when "000110111001000111" => data <= "000000";
				when "000110111001001000" => data <= "000000";
				when "000110111001001001" => data <= "000000";
				when "000110111001001010" => data <= "000000";
				when "000110111001001011" => data <= "000000";
				when "000110111001001100" => data <= "000000";
				when "000110111001001101" => data <= "000000";
				when "000110111001001110" => data <= "000000";
				when "000110111001001111" => data <= "000000";
				when "000110111001010000" => data <= "000000";
				when "000110111001010001" => data <= "000000";
				when "000110111001010010" => data <= "000000";
				when "000110111001010011" => data <= "000000";
				when "000110111001010100" => data <= "000000";
				when "000110111001010101" => data <= "000000";
				when "000110111001010110" => data <= "000000";
				when "000110111001010111" => data <= "000000";
				when "000110111001011000" => data <= "000000";
				when "000110111001011001" => data <= "000000";
				when "000110111001011010" => data <= "000000";
				when "000110111001011011" => data <= "000000";
				when "000110111001011100" => data <= "000000";
				when "000110111001011101" => data <= "000000";
				when "000110111001011110" => data <= "000000";
				when "000110111001011111" => data <= "000000";
				when "000110111001100000" => data <= "000000";
				when "000110111001100001" => data <= "000000";
				when "000110111001100010" => data <= "000000";
				when "000110111001100011" => data <= "000000";
				when "000110111001100100" => data <= "000000";
				when "000110111001100101" => data <= "000000";
				when "000110111001100110" => data <= "000000";
				when "000110111001100111" => data <= "000000";
				when "000110111001101000" => data <= "000000";
				when "000110111001101001" => data <= "000000";
				when "000110111001101010" => data <= "000000";
				when "000110111001101011" => data <= "000000";
				when "000110111001101100" => data <= "000000";
				when "000110111001101101" => data <= "000000";
				when "000110111001101110" => data <= "000000";
				when "000110111001101111" => data <= "000000";
				when "000110111001110000" => data <= "000000";
				when "000110111001110001" => data <= "000000";
				when "000110111001110010" => data <= "000000";
				when "000110111001110011" => data <= "000000";
				when "000110111001110100" => data <= "000000";
				when "000110111001110101" => data <= "000000";
				when "000110111001110110" => data <= "000000";
				when "000110111001110111" => data <= "000000";
				when "000110111001111000" => data <= "000000";
				when "000110111001111001" => data <= "000000";
				when "000110111001111010" => data <= "000000";
				when "000110111001111011" => data <= "000000";
				when "000110111001111100" => data <= "000000";
				when "000110111001111101" => data <= "000000";
				when "000110111001111110" => data <= "000000";
				when "000110111001111111" => data <= "000000";
				when "000110111010000000" => data <= "000000";
				when "000110111010000001" => data <= "000000";
				when "000110111010000010" => data <= "000000";
				when "000110111010000011" => data <= "000000";
				when "000110111010000100" => data <= "000000";
				when "000110111010000101" => data <= "000000";
				when "000110111010000110" => data <= "000000";
				when "000110111010000111" => data <= "000000";
				when "000110111010001000" => data <= "000000";
				when "000110111010001001" => data <= "000000";
				when "000110111010001010" => data <= "000000";
				when "000110111010001011" => data <= "000000";
				when "000110111010001100" => data <= "000000";
				when "000110111010001101" => data <= "000000";
				when "000110111010001110" => data <= "000000";
				when "000110111010001111" => data <= "000000";
				when "000110111010010000" => data <= "000000";
				when "000110111010010001" => data <= "000000";
				when "000110111010010010" => data <= "000000";
				when "000110111010010011" => data <= "000000";
				when "000110111010010100" => data <= "000000";
				when "000110111010010101" => data <= "000000";
				when "000110111010010110" => data <= "000000";
				when "000110111010010111" => data <= "000000";
				when "000110111010011000" => data <= "000000";
				when "000110111010011001" => data <= "000000";
				when "000110111010011010" => data <= "000000";
				when "000110111010011011" => data <= "000000";
				when "000110111010011100" => data <= "000000";
				when "000110111010011101" => data <= "000000";
				when "000110111010011110" => data <= "000000";
				when "000110111010011111" => data <= "000000";
				when "000111000000000000" => data <= "000000";
				when "000111000000000001" => data <= "000000";
				when "000111000000000010" => data <= "000000";
				when "000111000000000011" => data <= "000000";
				when "000111000000000100" => data <= "000000";
				when "000111000000000101" => data <= "000000";
				when "000111000000000110" => data <= "000000";
				when "000111000000000111" => data <= "000000";
				when "000111000000001000" => data <= "000000";
				when "000111000000001001" => data <= "000000";
				when "000111000000001010" => data <= "000000";
				when "000111000000001011" => data <= "000000";
				when "000111000000001100" => data <= "000000";
				when "000111000000001101" => data <= "000000";
				when "000111000000001110" => data <= "000000";
				when "000111000000001111" => data <= "000000";
				when "000111000000010000" => data <= "000000";
				when "000111000000010001" => data <= "000000";
				when "000111000000010010" => data <= "000000";
				when "000111000000010011" => data <= "000000";
				when "000111000000010100" => data <= "000000";
				when "000111000000010101" => data <= "000000";
				when "000111000000010110" => data <= "000000";
				when "000111000000010111" => data <= "000000";
				when "000111000000011000" => data <= "000000";
				when "000111000000011001" => data <= "000000";
				when "000111000000011010" => data <= "000000";
				when "000111000000011011" => data <= "000000";
				when "000111000000011100" => data <= "000000";
				when "000111000000011101" => data <= "000000";
				when "000111000000011110" => data <= "000000";
				when "000111000000011111" => data <= "000000";
				when "000111000000100000" => data <= "000000";
				when "000111000000100001" => data <= "000000";
				when "000111000000100010" => data <= "000000";
				when "000111000000100011" => data <= "000000";
				when "000111000000100100" => data <= "000000";
				when "000111000000100101" => data <= "000000";
				when "000111000000100110" => data <= "000000";
				when "000111000000100111" => data <= "000000";
				when "000111000000101000" => data <= "000000";
				when "000111000000101001" => data <= "000000";
				when "000111000000101010" => data <= "000000";
				when "000111000000101011" => data <= "000000";
				when "000111000000101100" => data <= "000000";
				when "000111000000101101" => data <= "000000";
				when "000111000000101110" => data <= "000000";
				when "000111000000101111" => data <= "000000";
				when "000111000000110000" => data <= "000000";
				when "000111000000110001" => data <= "000000";
				when "000111000000110010" => data <= "000000";
				when "000111000000110011" => data <= "000000";
				when "000111000000110100" => data <= "000000";
				when "000111000000110101" => data <= "000000";
				when "000111000000110110" => data <= "000000";
				when "000111000000110111" => data <= "000000";
				when "000111000000111000" => data <= "000000";
				when "000111000000111001" => data <= "000000";
				when "000111000000111010" => data <= "000000";
				when "000111000000111011" => data <= "000000";
				when "000111000000111100" => data <= "000000";
				when "000111000000111101" => data <= "000000";
				when "000111000000111110" => data <= "000000";
				when "000111000000111111" => data <= "000000";
				when "000111000001000000" => data <= "000000";
				when "000111000001000001" => data <= "000000";
				when "000111000001000010" => data <= "000000";
				when "000111000001000011" => data <= "000000";
				when "000111000001000100" => data <= "000000";
				when "000111000001000101" => data <= "000000";
				when "000111000001000110" => data <= "000000";
				when "000111000001000111" => data <= "000000";
				when "000111000001001000" => data <= "000000";
				when "000111000001001001" => data <= "000000";
				when "000111000001001010" => data <= "000000";
				when "000111000001001011" => data <= "000000";
				when "000111000001001100" => data <= "000000";
				when "000111000001001101" => data <= "000000";
				when "000111000001001110" => data <= "000000";
				when "000111000001001111" => data <= "000000";
				when "000111000001010000" => data <= "000000";
				when "000111000001010001" => data <= "000000";
				when "000111000001010010" => data <= "000000";
				when "000111000001010011" => data <= "000000";
				when "000111000001010100" => data <= "000000";
				when "000111000001010101" => data <= "000000";
				when "000111000001010110" => data <= "000000";
				when "000111000001010111" => data <= "000000";
				when "000111000001011000" => data <= "000000";
				when "000111000001011001" => data <= "000000";
				when "000111000001011010" => data <= "000000";
				when "000111000001011011" => data <= "000000";
				when "000111000001011100" => data <= "000000";
				when "000111000001011101" => data <= "000000";
				when "000111000001011110" => data <= "000000";
				when "000111000001011111" => data <= "000000";
				when "000111000001100000" => data <= "000000";
				when "000111000001100001" => data <= "000000";
				when "000111000001100010" => data <= "000000";
				when "000111000001100011" => data <= "000000";
				when "000111000001100100" => data <= "000000";
				when "000111000001100101" => data <= "000000";
				when "000111000001100110" => data <= "000000";
				when "000111000001100111" => data <= "000000";
				when "000111000001101000" => data <= "000000";
				when "000111000001101001" => data <= "000000";
				when "000111000001101010" => data <= "000000";
				when "000111000001101011" => data <= "000000";
				when "000111000001101100" => data <= "000000";
				when "000111000001101101" => data <= "000000";
				when "000111000001101110" => data <= "000000";
				when "000111000001101111" => data <= "000000";
				when "000111000001110000" => data <= "000000";
				when "000111000001110001" => data <= "000000";
				when "000111000001110010" => data <= "000000";
				when "000111000001110011" => data <= "000000";
				when "000111000001110100" => data <= "000000";
				when "000111000001110101" => data <= "000000";
				when "000111000001110110" => data <= "000000";
				when "000111000001110111" => data <= "000000";
				when "000111000001111000" => data <= "000000";
				when "000111000001111001" => data <= "000000";
				when "000111000001111010" => data <= "000000";
				when "000111000001111011" => data <= "000000";
				when "000111000001111100" => data <= "000000";
				when "000111000001111101" => data <= "000000";
				when "000111000001111110" => data <= "000000";
				when "000111000001111111" => data <= "000000";
				when "000111000010000000" => data <= "000000";
				when "000111000010000001" => data <= "000000";
				when "000111000010000010" => data <= "000000";
				when "000111000010000011" => data <= "000000";
				when "000111000010000100" => data <= "000000";
				when "000111000010000101" => data <= "000000";
				when "000111000010000110" => data <= "000000";
				when "000111000010000111" => data <= "000000";
				when "000111000010001000" => data <= "000000";
				when "000111000010001001" => data <= "000000";
				when "000111000010001010" => data <= "000000";
				when "000111000010001011" => data <= "000000";
				when "000111000010001100" => data <= "000000";
				when "000111000010001101" => data <= "000000";
				when "000111000010001110" => data <= "000000";
				when "000111000010001111" => data <= "000000";
				when "000111000010010000" => data <= "000000";
				when "000111000010010001" => data <= "000000";
				when "000111000010010010" => data <= "000000";
				when "000111000010010011" => data <= "000000";
				when "000111000010010100" => data <= "000000";
				when "000111000010010101" => data <= "000000";
				when "000111000010010110" => data <= "000000";
				when "000111000010010111" => data <= "000000";
				when "000111000010011000" => data <= "000000";
				when "000111000010011001" => data <= "000000";
				when "000111000010011010" => data <= "000000";
				when "000111000010011011" => data <= "000000";
				when "000111000010011100" => data <= "000000";
				when "000111000010011101" => data <= "000000";
				when "000111000010011110" => data <= "000000";
				when "000111000010011111" => data <= "000000";
				when "000111001000000000" => data <= "000000";
				when "000111001000000001" => data <= "000000";
				when "000111001000000010" => data <= "000000";
				when "000111001000000011" => data <= "000000";
				when "000111001000000100" => data <= "000000";
				when "000111001000000101" => data <= "000000";
				when "000111001000000110" => data <= "000000";
				when "000111001000000111" => data <= "000000";
				when "000111001000001000" => data <= "000000";
				when "000111001000001001" => data <= "000000";
				when "000111001000001010" => data <= "000000";
				when "000111001000001011" => data <= "000000";
				when "000111001000001100" => data <= "000000";
				when "000111001000001101" => data <= "000000";
				when "000111001000001110" => data <= "000000";
				when "000111001000001111" => data <= "000000";
				when "000111001000010000" => data <= "000000";
				when "000111001000010001" => data <= "000000";
				when "000111001000010010" => data <= "000000";
				when "000111001000010011" => data <= "000000";
				when "000111001000010100" => data <= "000000";
				when "000111001000010101" => data <= "000000";
				when "000111001000010110" => data <= "000000";
				when "000111001000010111" => data <= "000000";
				when "000111001000011000" => data <= "000000";
				when "000111001000011001" => data <= "000000";
				when "000111001000011010" => data <= "000000";
				when "000111001000011011" => data <= "000000";
				when "000111001000011100" => data <= "000000";
				when "000111001000011101" => data <= "000000";
				when "000111001000011110" => data <= "000000";
				when "000111001000011111" => data <= "000000";
				when "000111001000100000" => data <= "000000";
				when "000111001000100001" => data <= "000000";
				when "000111001000100010" => data <= "000000";
				when "000111001000100011" => data <= "000000";
				when "000111001000100100" => data <= "000000";
				when "000111001000100101" => data <= "000000";
				when "000111001000100110" => data <= "000000";
				when "000111001000100111" => data <= "000000";
				when "000111001000101000" => data <= "000000";
				when "000111001000101001" => data <= "000000";
				when "000111001000101010" => data <= "000000";
				when "000111001000101011" => data <= "000000";
				when "000111001000101100" => data <= "000000";
				when "000111001000101101" => data <= "000000";
				when "000111001000101110" => data <= "000000";
				when "000111001000101111" => data <= "000000";
				when "000111001000110000" => data <= "000000";
				when "000111001000110001" => data <= "000000";
				when "000111001000110010" => data <= "000000";
				when "000111001000110011" => data <= "000000";
				when "000111001000110100" => data <= "000000";
				when "000111001000110101" => data <= "000000";
				when "000111001000110110" => data <= "000000";
				when "000111001000110111" => data <= "000000";
				when "000111001000111000" => data <= "000000";
				when "000111001000111001" => data <= "000000";
				when "000111001000111010" => data <= "000000";
				when "000111001000111011" => data <= "000000";
				when "000111001000111100" => data <= "000000";
				when "000111001000111101" => data <= "000000";
				when "000111001000111110" => data <= "000000";
				when "000111001000111111" => data <= "000000";
				when "000111001001000000" => data <= "000000";
				when "000111001001000001" => data <= "000000";
				when "000111001001000010" => data <= "000000";
				when "000111001001000011" => data <= "000000";
				when "000111001001000100" => data <= "000000";
				when "000111001001000101" => data <= "000000";
				when "000111001001000110" => data <= "000000";
				when "000111001001000111" => data <= "000000";
				when "000111001001001000" => data <= "000000";
				when "000111001001001001" => data <= "000000";
				when "000111001001001010" => data <= "000000";
				when "000111001001001011" => data <= "000000";
				when "000111001001001100" => data <= "000000";
				when "000111001001001101" => data <= "000000";
				when "000111001001001110" => data <= "000000";
				when "000111001001001111" => data <= "000000";
				when "000111001001010000" => data <= "000000";
				when "000111001001010001" => data <= "000000";
				when "000111001001010010" => data <= "000000";
				when "000111001001010011" => data <= "000000";
				when "000111001001010100" => data <= "000000";
				when "000111001001010101" => data <= "000000";
				when "000111001001010110" => data <= "000000";
				when "000111001001010111" => data <= "000000";
				when "000111001001011000" => data <= "000000";
				when "000111001001011001" => data <= "000000";
				when "000111001001011010" => data <= "000000";
				when "000111001001011011" => data <= "000000";
				when "000111001001011100" => data <= "000000";
				when "000111001001011101" => data <= "000000";
				when "000111001001011110" => data <= "000000";
				when "000111001001011111" => data <= "000000";
				when "000111001001100000" => data <= "000000";
				when "000111001001100001" => data <= "000000";
				when "000111001001100010" => data <= "000000";
				when "000111001001100011" => data <= "000000";
				when "000111001001100100" => data <= "000000";
				when "000111001001100101" => data <= "000000";
				when "000111001001100110" => data <= "000000";
				when "000111001001100111" => data <= "000000";
				when "000111001001101000" => data <= "000000";
				when "000111001001101001" => data <= "000000";
				when "000111001001101010" => data <= "000000";
				when "000111001001101011" => data <= "000000";
				when "000111001001101100" => data <= "000000";
				when "000111001001101101" => data <= "000000";
				when "000111001001101110" => data <= "000000";
				when "000111001001101111" => data <= "000000";
				when "000111001001110000" => data <= "000000";
				when "000111001001110001" => data <= "000000";
				when "000111001001110010" => data <= "000000";
				when "000111001001110011" => data <= "000000";
				when "000111001001110100" => data <= "000000";
				when "000111001001110101" => data <= "000000";
				when "000111001001110110" => data <= "000000";
				when "000111001001110111" => data <= "000000";
				when "000111001001111000" => data <= "000000";
				when "000111001001111001" => data <= "000000";
				when "000111001001111010" => data <= "000000";
				when "000111001001111011" => data <= "000000";
				when "000111001001111100" => data <= "000000";
				when "000111001001111101" => data <= "000000";
				when "000111001001111110" => data <= "000000";
				when "000111001001111111" => data <= "000000";
				when "000111001010000000" => data <= "000000";
				when "000111001010000001" => data <= "000000";
				when "000111001010000010" => data <= "000000";
				when "000111001010000011" => data <= "000000";
				when "000111001010000100" => data <= "000000";
				when "000111001010000101" => data <= "000000";
				when "000111001010000110" => data <= "000000";
				when "000111001010000111" => data <= "000000";
				when "000111001010001000" => data <= "000000";
				when "000111001010001001" => data <= "000000";
				when "000111001010001010" => data <= "000000";
				when "000111001010001011" => data <= "000000";
				when "000111001010001100" => data <= "000000";
				when "000111001010001101" => data <= "000000";
				when "000111001010001110" => data <= "000000";
				when "000111001010001111" => data <= "000000";
				when "000111001010010000" => data <= "000000";
				when "000111001010010001" => data <= "000000";
				when "000111001010010010" => data <= "000000";
				when "000111001010010011" => data <= "000000";
				when "000111001010010100" => data <= "000000";
				when "000111001010010101" => data <= "000000";
				when "000111001010010110" => data <= "000000";
				when "000111001010010111" => data <= "000000";
				when "000111001010011000" => data <= "000000";
				when "000111001010011001" => data <= "000000";
				when "000111001010011010" => data <= "000000";
				when "000111001010011011" => data <= "000000";
				when "000111001010011100" => data <= "000000";
				when "000111001010011101" => data <= "000000";
				when "000111001010011110" => data <= "000000";
				when "000111001010011111" => data <= "000000";
				when "000111010000000000" => data <= "000000";
				when "000111010000000001" => data <= "000000";
				when "000111010000000010" => data <= "000000";
				when "000111010000000011" => data <= "000000";
				when "000111010000000100" => data <= "000000";
				when "000111010000000101" => data <= "000000";
				when "000111010000000110" => data <= "000000";
				when "000111010000000111" => data <= "000000";
				when "000111010000001000" => data <= "000000";
				when "000111010000001001" => data <= "000000";
				when "000111010000001010" => data <= "000000";
				when "000111010000001011" => data <= "000000";
				when "000111010000001100" => data <= "000000";
				when "000111010000001101" => data <= "000000";
				when "000111010000001110" => data <= "000000";
				when "000111010000001111" => data <= "000000";
				when "000111010000010000" => data <= "000000";
				when "000111010000010001" => data <= "000000";
				when "000111010000010010" => data <= "000000";
				when "000111010000010011" => data <= "000000";
				when "000111010000010100" => data <= "000000";
				when "000111010000010101" => data <= "000000";
				when "000111010000010110" => data <= "000000";
				when "000111010000010111" => data <= "000000";
				when "000111010000011000" => data <= "000000";
				when "000111010000011001" => data <= "000000";
				when "000111010000011010" => data <= "000000";
				when "000111010000011011" => data <= "000000";
				when "000111010000011100" => data <= "000000";
				when "000111010000011101" => data <= "000000";
				when "000111010000011110" => data <= "000000";
				when "000111010000011111" => data <= "000000";
				when "000111010000100000" => data <= "000000";
				when "000111010000100001" => data <= "000000";
				when "000111010000100010" => data <= "000000";
				when "000111010000100011" => data <= "000000";
				when "000111010000100100" => data <= "000000";
				when "000111010000100101" => data <= "000000";
				when "000111010000100110" => data <= "000000";
				when "000111010000100111" => data <= "000000";
				when "000111010000101000" => data <= "000000";
				when "000111010000101001" => data <= "000000";
				when "000111010000101010" => data <= "000000";
				when "000111010000101011" => data <= "000000";
				when "000111010000101100" => data <= "000000";
				when "000111010000101101" => data <= "000000";
				when "000111010000101110" => data <= "000000";
				when "000111010000101111" => data <= "000000";
				when "000111010000110000" => data <= "000000";
				when "000111010000110001" => data <= "000000";
				when "000111010000110010" => data <= "000000";
				when "000111010000110011" => data <= "000000";
				when "000111010000110100" => data <= "000000";
				when "000111010000110101" => data <= "000000";
				when "000111010000110110" => data <= "000000";
				when "000111010000110111" => data <= "000000";
				when "000111010000111000" => data <= "000000";
				when "000111010000111001" => data <= "000000";
				when "000111010000111010" => data <= "000000";
				when "000111010000111011" => data <= "000000";
				when "000111010000111100" => data <= "000000";
				when "000111010000111101" => data <= "000000";
				when "000111010000111110" => data <= "000000";
				when "000111010000111111" => data <= "000000";
				when "000111010001000000" => data <= "000000";
				when "000111010001000001" => data <= "000000";
				when "000111010001000010" => data <= "000000";
				when "000111010001000011" => data <= "000000";
				when "000111010001000100" => data <= "000000";
				when "000111010001000101" => data <= "000000";
				when "000111010001000110" => data <= "000000";
				when "000111010001000111" => data <= "000000";
				when "000111010001001000" => data <= "000000";
				when "000111010001001001" => data <= "000000";
				when "000111010001001010" => data <= "000000";
				when "000111010001001011" => data <= "000000";
				when "000111010001001100" => data <= "000000";
				when "000111010001001101" => data <= "000000";
				when "000111010001001110" => data <= "000000";
				when "000111010001001111" => data <= "000000";
				when "000111010001010000" => data <= "000000";
				when "000111010001010001" => data <= "000000";
				when "000111010001010010" => data <= "000000";
				when "000111010001010011" => data <= "000000";
				when "000111010001010100" => data <= "000000";
				when "000111010001010101" => data <= "000000";
				when "000111010001010110" => data <= "000000";
				when "000111010001010111" => data <= "000000";
				when "000111010001011000" => data <= "000000";
				when "000111010001011001" => data <= "000000";
				when "000111010001011010" => data <= "000000";
				when "000111010001011011" => data <= "000000";
				when "000111010001011100" => data <= "000000";
				when "000111010001011101" => data <= "000000";
				when "000111010001011110" => data <= "000000";
				when "000111010001011111" => data <= "000000";
				when "000111010001100000" => data <= "000000";
				when "000111010001100001" => data <= "000000";
				when "000111010001100010" => data <= "000000";
				when "000111010001100011" => data <= "000000";
				when "000111010001100100" => data <= "000000";
				when "000111010001100101" => data <= "000000";
				when "000111010001100110" => data <= "000000";
				when "000111010001100111" => data <= "000000";
				when "000111010001101000" => data <= "000000";
				when "000111010001101001" => data <= "000000";
				when "000111010001101010" => data <= "000000";
				when "000111010001101011" => data <= "000000";
				when "000111010001101100" => data <= "000000";
				when "000111010001101101" => data <= "000000";
				when "000111010001101110" => data <= "000000";
				when "000111010001101111" => data <= "000000";
				when "000111010001110000" => data <= "000000";
				when "000111010001110001" => data <= "000000";
				when "000111010001110010" => data <= "000000";
				when "000111010001110011" => data <= "000000";
				when "000111010001110100" => data <= "000000";
				when "000111010001110101" => data <= "000000";
				when "000111010001110110" => data <= "000000";
				when "000111010001110111" => data <= "000000";
				when "000111010001111000" => data <= "000000";
				when "000111010001111001" => data <= "000000";
				when "000111010001111010" => data <= "000000";
				when "000111010001111011" => data <= "000000";
				when "000111010001111100" => data <= "000000";
				when "000111010001111101" => data <= "000000";
				when "000111010001111110" => data <= "000000";
				when "000111010001111111" => data <= "000000";
				when "000111010010000000" => data <= "000000";
				when "000111010010000001" => data <= "000000";
				when "000111010010000010" => data <= "000000";
				when "000111010010000011" => data <= "000000";
				when "000111010010000100" => data <= "000000";
				when "000111010010000101" => data <= "000000";
				when "000111010010000110" => data <= "000000";
				when "000111010010000111" => data <= "000000";
				when "000111010010001000" => data <= "000000";
				when "000111010010001001" => data <= "000000";
				when "000111010010001010" => data <= "000000";
				when "000111010010001011" => data <= "000000";
				when "000111010010001100" => data <= "000000";
				when "000111010010001101" => data <= "000000";
				when "000111010010001110" => data <= "000000";
				when "000111010010001111" => data <= "000000";
				when "000111010010010000" => data <= "000000";
				when "000111010010010001" => data <= "000000";
				when "000111010010010010" => data <= "000000";
				when "000111010010010011" => data <= "000000";
				when "000111010010010100" => data <= "000000";
				when "000111010010010101" => data <= "000000";
				when "000111010010010110" => data <= "000000";
				when "000111010010010111" => data <= "000000";
				when "000111010010011000" => data <= "000000";
				when "000111010010011001" => data <= "000000";
				when "000111010010011010" => data <= "000000";
				when "000111010010011011" => data <= "000000";
				when "000111010010011100" => data <= "000000";
				when "000111010010011101" => data <= "000000";
				when "000111010010011110" => data <= "000000";
				when "000111010010011111" => data <= "000000";
				when "000111011000000000" => data <= "000000";
				when "000111011000000001" => data <= "000000";
				when "000111011000000010" => data <= "000000";
				when "000111011000000011" => data <= "000000";
				when "000111011000000100" => data <= "000000";
				when "000111011000000101" => data <= "000000";
				when "000111011000000110" => data <= "000000";
				when "000111011000000111" => data <= "000000";
				when "000111011000001000" => data <= "000000";
				when "000111011000001001" => data <= "000000";
				when "000111011000001010" => data <= "000000";
				when "000111011000001011" => data <= "000000";
				when "000111011000001100" => data <= "000000";
				when "000111011000001101" => data <= "000000";
				when "000111011000001110" => data <= "000000";
				when "000111011000001111" => data <= "000000";
				when "000111011000010000" => data <= "000000";
				when "000111011000010001" => data <= "000000";
				when "000111011000010010" => data <= "000000";
				when "000111011000010011" => data <= "000000";
				when "000111011000010100" => data <= "000000";
				when "000111011000010101" => data <= "000000";
				when "000111011000010110" => data <= "000000";
				when "000111011000010111" => data <= "000000";
				when "000111011000011000" => data <= "000000";
				when "000111011000011001" => data <= "000000";
				when "000111011000011010" => data <= "000000";
				when "000111011000011011" => data <= "000000";
				when "000111011000011100" => data <= "000000";
				when "000111011000011101" => data <= "000000";
				when "000111011000011110" => data <= "000000";
				when "000111011000011111" => data <= "000000";
				when "000111011000100000" => data <= "000000";
				when "000111011000100001" => data <= "000000";
				when "000111011000100010" => data <= "000000";
				when "000111011000100011" => data <= "000000";
				when "000111011000100100" => data <= "000000";
				when "000111011000100101" => data <= "000000";
				when "000111011000100110" => data <= "000000";
				when "000111011000100111" => data <= "000000";
				when "000111011000101000" => data <= "000000";
				when "000111011000101001" => data <= "000000";
				when "000111011000101010" => data <= "000000";
				when "000111011000101011" => data <= "000000";
				when "000111011000101100" => data <= "000000";
				when "000111011000101101" => data <= "000000";
				when "000111011000101110" => data <= "000000";
				when "000111011000101111" => data <= "000000";
				when "000111011000110000" => data <= "000000";
				when "000111011000110001" => data <= "000000";
				when "000111011000110010" => data <= "000000";
				when "000111011000110011" => data <= "000000";
				when "000111011000110100" => data <= "000000";
				when "000111011000110101" => data <= "000000";
				when "000111011000110110" => data <= "000000";
				when "000111011000110111" => data <= "000000";
				when "000111011000111000" => data <= "000000";
				when "000111011000111001" => data <= "000000";
				when "000111011000111010" => data <= "000000";
				when "000111011000111011" => data <= "000000";
				when "000111011000111100" => data <= "000000";
				when "000111011000111101" => data <= "000000";
				when "000111011000111110" => data <= "000000";
				when "000111011000111111" => data <= "000000";
				when "000111011001000000" => data <= "000000";
				when "000111011001000001" => data <= "000000";
				when "000111011001000010" => data <= "000000";
				when "000111011001000011" => data <= "000000";
				when "000111011001000100" => data <= "000000";
				when "000111011001000101" => data <= "000000";
				when "000111011001000110" => data <= "000000";
				when "000111011001000111" => data <= "000000";
				when "000111011001001000" => data <= "000000";
				when "000111011001001001" => data <= "000000";
				when "000111011001001010" => data <= "000000";
				when "000111011001001011" => data <= "000000";
				when "000111011001001100" => data <= "000000";
				when "000111011001001101" => data <= "000000";
				when "000111011001001110" => data <= "000000";
				when "000111011001001111" => data <= "000000";
				when "000111011001010000" => data <= "000000";
				when "000111011001010001" => data <= "000000";
				when "000111011001010010" => data <= "000000";
				when "000111011001010011" => data <= "000000";
				when "000111011001010100" => data <= "000000";
				when "000111011001010101" => data <= "000000";
				when "000111011001010110" => data <= "000000";
				when "000111011001010111" => data <= "000000";
				when "000111011001011000" => data <= "000000";
				when "000111011001011001" => data <= "000000";
				when "000111011001011010" => data <= "000000";
				when "000111011001011011" => data <= "000000";
				when "000111011001011100" => data <= "000000";
				when "000111011001011101" => data <= "000000";
				when "000111011001011110" => data <= "000000";
				when "000111011001011111" => data <= "000000";
				when "000111011001100000" => data <= "000000";
				when "000111011001100001" => data <= "000000";
				when "000111011001100010" => data <= "000000";
				when "000111011001100011" => data <= "000000";
				when "000111011001100100" => data <= "000000";
				when "000111011001100101" => data <= "000000";
				when "000111011001100110" => data <= "000000";
				when "000111011001100111" => data <= "000000";
				when "000111011001101000" => data <= "000000";
				when "000111011001101001" => data <= "000000";
				when "000111011001101010" => data <= "000000";
				when "000111011001101011" => data <= "000000";
				when "000111011001101100" => data <= "000000";
				when "000111011001101101" => data <= "000000";
				when "000111011001101110" => data <= "000000";
				when "000111011001101111" => data <= "000000";
				when "000111011001110000" => data <= "000000";
				when "000111011001110001" => data <= "000000";
				when "000111011001110010" => data <= "000000";
				when "000111011001110011" => data <= "000000";
				when "000111011001110100" => data <= "000000";
				when "000111011001110101" => data <= "000000";
				when "000111011001110110" => data <= "000000";
				when "000111011001110111" => data <= "000000";
				when "000111011001111000" => data <= "000000";
				when "000111011001111001" => data <= "000000";
				when "000111011001111010" => data <= "000000";
				when "000111011001111011" => data <= "000000";
				when "000111011001111100" => data <= "000000";
				when "000111011001111101" => data <= "000000";
				when "000111011001111110" => data <= "000000";
				when "000111011001111111" => data <= "000000";
				when "000111011010000000" => data <= "000000";
				when "000111011010000001" => data <= "000000";
				when "000111011010000010" => data <= "000000";
				when "000111011010000011" => data <= "000000";
				when "000111011010000100" => data <= "000000";
				when "000111011010000101" => data <= "000000";
				when "000111011010000110" => data <= "000000";
				when "000111011010000111" => data <= "000000";
				when "000111011010001000" => data <= "000000";
				when "000111011010001001" => data <= "000000";
				when "000111011010001010" => data <= "000000";
				when "000111011010001011" => data <= "000000";
				when "000111011010001100" => data <= "000000";
				when "000111011010001101" => data <= "000000";
				when "000111011010001110" => data <= "000000";
				when "000111011010001111" => data <= "000000";
				when "000111011010010000" => data <= "000000";
				when "000111011010010001" => data <= "000000";
				when "000111011010010010" => data <= "000000";
				when "000111011010010011" => data <= "000000";
				when "000111011010010100" => data <= "000000";
				when "000111011010010101" => data <= "000000";
				when "000111011010010110" => data <= "000000";
				when "000111011010010111" => data <= "000000";
				when "000111011010011000" => data <= "000000";
				when "000111011010011001" => data <= "000000";
				when "000111011010011010" => data <= "000000";
				when "000111011010011011" => data <= "000000";
				when "000111011010011100" => data <= "000000";
				when "000111011010011101" => data <= "000000";
				when "000111011010011110" => data <= "000000";
				when "000111011010011111" => data <= "000000";
				when "000111100000000000" => data <= "000000";
				when "000111100000000001" => data <= "000000";
				when "000111100000000010" => data <= "000000";
				when "000111100000000011" => data <= "000000";
				when "000111100000000100" => data <= "000000";
				when "000111100000000101" => data <= "000000";
				when "000111100000000110" => data <= "000000";
				when "000111100000000111" => data <= "000000";
				when "000111100000001000" => data <= "000000";
				when "000111100000001001" => data <= "000000";
				when "000111100000001010" => data <= "000000";
				when "000111100000001011" => data <= "000000";
				when "000111100000001100" => data <= "000000";
				when "000111100000001101" => data <= "000000";
				when "000111100000001110" => data <= "000000";
				when "000111100000001111" => data <= "000000";
				when "000111100000010000" => data <= "000000";
				when "000111100000010001" => data <= "000000";
				when "000111100000010010" => data <= "000000";
				when "000111100000010011" => data <= "000000";
				when "000111100000010100" => data <= "000000";
				when "000111100000010101" => data <= "000000";
				when "000111100000010110" => data <= "000000";
				when "000111100000010111" => data <= "000000";
				when "000111100000011000" => data <= "000000";
				when "000111100000011001" => data <= "000000";
				when "000111100000011010" => data <= "000000";
				when "000111100000011011" => data <= "000000";
				when "000111100000011100" => data <= "000000";
				when "000111100000011101" => data <= "000000";
				when "000111100000011110" => data <= "000000";
				when "000111100000011111" => data <= "000000";
				when "000111100000100000" => data <= "000000";
				when "000111100000100001" => data <= "000000";
				when "000111100000100010" => data <= "000000";
				when "000111100000100011" => data <= "000000";
				when "000111100000100100" => data <= "000000";
				when "000111100000100101" => data <= "000000";
				when "000111100000100110" => data <= "000000";
				when "000111100000100111" => data <= "000000";
				when "000111100000101000" => data <= "000000";
				when "000111100000101001" => data <= "000000";
				when "000111100000101010" => data <= "000000";
				when "000111100000101011" => data <= "000000";
				when "000111100000101100" => data <= "000000";
				when "000111100000101101" => data <= "000000";
				when "000111100000101110" => data <= "000000";
				when "000111100000101111" => data <= "000000";
				when "000111100000110000" => data <= "000000";
				when "000111100000110001" => data <= "000000";
				when "000111100000110010" => data <= "000000";
				when "000111100000110011" => data <= "000000";
				when "000111100000110100" => data <= "000000";
				when "000111100000110101" => data <= "000000";
				when "000111100000110110" => data <= "000000";
				when "000111100000110111" => data <= "000000";
				when "000111100000111000" => data <= "000000";
				when "000111100000111001" => data <= "000000";
				when "000111100000111010" => data <= "000000";
				when "000111100000111011" => data <= "000000";
				when "000111100000111100" => data <= "000000";
				when "000111100000111101" => data <= "000000";
				when "000111100000111110" => data <= "000000";
				when "000111100000111111" => data <= "000000";
				when "000111100001000000" => data <= "000000";
				when "000111100001000001" => data <= "000000";
				when "000111100001000010" => data <= "000000";
				when "000111100001000011" => data <= "000000";
				when "000111100001000100" => data <= "000000";
				when "000111100001000101" => data <= "000000";
				when "000111100001000110" => data <= "000000";
				when "000111100001000111" => data <= "000000";
				when "000111100001001000" => data <= "000000";
				when "000111100001001001" => data <= "000000";
				when "000111100001001010" => data <= "000000";
				when "000111100001001011" => data <= "000000";
				when "000111100001001100" => data <= "000000";
				when "000111100001001101" => data <= "000000";
				when "000111100001001110" => data <= "000000";
				when "000111100001001111" => data <= "000000";
				when "000111100001010000" => data <= "000000";
				when "000111100001010001" => data <= "000000";
				when "000111100001010010" => data <= "000000";
				when "000111100001010011" => data <= "000000";
				when "000111100001010100" => data <= "000000";
				when "000111100001010101" => data <= "000000";
				when "000111100001010110" => data <= "000000";
				when "000111100001010111" => data <= "000000";
				when "000111100001011000" => data <= "000000";
				when "000111100001011001" => data <= "000000";
				when "000111100001011010" => data <= "000000";
				when "000111100001011011" => data <= "000000";
				when "000111100001011100" => data <= "000000";
				when "000111100001011101" => data <= "000000";
				when "000111100001011110" => data <= "000000";
				when "000111100001011111" => data <= "000000";
				when "000111100001100000" => data <= "000000";
				when "000111100001100001" => data <= "000000";
				when "000111100001100010" => data <= "000000";
				when "000111100001100011" => data <= "000000";
				when "000111100001100100" => data <= "000000";
				when "000111100001100101" => data <= "000000";
				when "000111100001100110" => data <= "000000";
				when "000111100001100111" => data <= "000000";
				when "000111100001101000" => data <= "000000";
				when "000111100001101001" => data <= "000000";
				when "000111100001101010" => data <= "000000";
				when "000111100001101011" => data <= "000000";
				when "000111100001101100" => data <= "000000";
				when "000111100001101101" => data <= "000000";
				when "000111100001101110" => data <= "000000";
				when "000111100001101111" => data <= "000000";
				when "000111100001110000" => data <= "000000";
				when "000111100001110001" => data <= "000000";
				when "000111100001110010" => data <= "000000";
				when "000111100001110011" => data <= "000000";
				when "000111100001110100" => data <= "000000";
				when "000111100001110101" => data <= "000000";
				when "000111100001110110" => data <= "000000";
				when "000111100001110111" => data <= "000000";
				when "000111100001111000" => data <= "000000";
				when "000111100001111001" => data <= "000000";
				when "000111100001111010" => data <= "000000";
				when "000111100001111011" => data <= "000000";
				when "000111100001111100" => data <= "000000";
				when "000111100001111101" => data <= "000000";
				when "000111100001111110" => data <= "000000";
				when "000111100001111111" => data <= "000000";
				when "000111100010000000" => data <= "000000";
				when "000111100010000001" => data <= "000000";
				when "000111100010000010" => data <= "000000";
				when "000111100010000011" => data <= "000000";
				when "000111100010000100" => data <= "000000";
				when "000111100010000101" => data <= "000000";
				when "000111100010000110" => data <= "000000";
				when "000111100010000111" => data <= "000000";
				when "000111100010001000" => data <= "000000";
				when "000111100010001001" => data <= "000000";
				when "000111100010001010" => data <= "000000";
				when "000111100010001011" => data <= "000000";
				when "000111100010001100" => data <= "000000";
				when "000111100010001101" => data <= "000000";
				when "000111100010001110" => data <= "000000";
				when "000111100010001111" => data <= "000000";
				when "000111100010010000" => data <= "000000";
				when "000111100010010001" => data <= "000000";
				when "000111100010010010" => data <= "000000";
				when "000111100010010011" => data <= "000000";
				when "000111100010010100" => data <= "000000";
				when "000111100010010101" => data <= "000000";
				when "000111100010010110" => data <= "000000";
				when "000111100010010111" => data <= "000000";
				when "000111100010011000" => data <= "000000";
				when "000111100010011001" => data <= "000000";
				when "000111100010011010" => data <= "000000";
				when "000111100010011011" => data <= "000000";
				when "000111100010011100" => data <= "000000";
				when "000111100010011101" => data <= "000000";
				when "000111100010011110" => data <= "000000";
				when "000111100010011111" => data <= "000000";
				when "000111101000000000" => data <= "000000";
				when "000111101000000001" => data <= "000000";
				when "000111101000000010" => data <= "000000";
				when "000111101000000011" => data <= "000000";
				when "000111101000000100" => data <= "000000";
				when "000111101000000101" => data <= "000000";
				when "000111101000000110" => data <= "000000";
				when "000111101000000111" => data <= "000000";
				when "000111101000001000" => data <= "000000";
				when "000111101000001001" => data <= "000000";
				when "000111101000001010" => data <= "000000";
				when "000111101000001011" => data <= "000000";
				when "000111101000001100" => data <= "000000";
				when "000111101000001101" => data <= "000000";
				when "000111101000001110" => data <= "000000";
				when "000111101000001111" => data <= "000000";
				when "000111101000010000" => data <= "000000";
				when "000111101000010001" => data <= "000000";
				when "000111101000010010" => data <= "000000";
				when "000111101000010011" => data <= "000000";
				when "000111101000010100" => data <= "000000";
				when "000111101000010101" => data <= "000000";
				when "000111101000010110" => data <= "000000";
				when "000111101000010111" => data <= "000000";
				when "000111101000011000" => data <= "000000";
				when "000111101000011001" => data <= "000000";
				when "000111101000011010" => data <= "000000";
				when "000111101000011011" => data <= "000000";
				when "000111101000011100" => data <= "000000";
				when "000111101000011101" => data <= "000000";
				when "000111101000011110" => data <= "000000";
				when "000111101000011111" => data <= "000000";
				when "000111101000100000" => data <= "000000";
				when "000111101000100001" => data <= "000000";
				when "000111101000100010" => data <= "000000";
				when "000111101000100011" => data <= "000000";
				when "000111101000100100" => data <= "000000";
				when "000111101000100101" => data <= "000000";
				when "000111101000100110" => data <= "000000";
				when "000111101000100111" => data <= "000000";
				when "000111101000101000" => data <= "000000";
				when "000111101000101001" => data <= "000000";
				when "000111101000101010" => data <= "000000";
				when "000111101000101011" => data <= "000000";
				when "000111101000101100" => data <= "000000";
				when "000111101000101101" => data <= "000000";
				when "000111101000101110" => data <= "000000";
				when "000111101000101111" => data <= "000000";
				when "000111101000110000" => data <= "000000";
				when "000111101000110001" => data <= "000000";
				when "000111101000110010" => data <= "000000";
				when "000111101000110011" => data <= "000000";
				when "000111101000110100" => data <= "000000";
				when "000111101000110101" => data <= "000000";
				when "000111101000110110" => data <= "000000";
				when "000111101000110111" => data <= "000000";
				when "000111101000111000" => data <= "000000";
				when "000111101000111001" => data <= "000000";
				when "000111101000111010" => data <= "000000";
				when "000111101000111011" => data <= "000000";
				when "000111101000111100" => data <= "000000";
				when "000111101000111101" => data <= "000000";
				when "000111101000111110" => data <= "000000";
				when "000111101000111111" => data <= "000000";
				when "000111101001000000" => data <= "000000";
				when "000111101001000001" => data <= "000000";
				when "000111101001000010" => data <= "000000";
				when "000111101001000011" => data <= "000000";
				when "000111101001000100" => data <= "000000";
				when "000111101001000101" => data <= "000000";
				when "000111101001000110" => data <= "000000";
				when "000111101001000111" => data <= "000000";
				when "000111101001001000" => data <= "000000";
				when "000111101001001001" => data <= "000000";
				when "000111101001001010" => data <= "000000";
				when "000111101001001011" => data <= "000000";
				when "000111101001001100" => data <= "000000";
				when "000111101001001101" => data <= "000000";
				when "000111101001001110" => data <= "000000";
				when "000111101001001111" => data <= "000000";
				when "000111101001010000" => data <= "000000";
				when "000111101001010001" => data <= "000000";
				when "000111101001010010" => data <= "000000";
				when "000111101001010011" => data <= "000000";
				when "000111101001010100" => data <= "000000";
				when "000111101001010101" => data <= "000000";
				when "000111101001010110" => data <= "000000";
				when "000111101001010111" => data <= "000000";
				when "000111101001011000" => data <= "000000";
				when "000111101001011001" => data <= "000000";
				when "000111101001011010" => data <= "000000";
				when "000111101001011011" => data <= "000000";
				when "000111101001011100" => data <= "000000";
				when "000111101001011101" => data <= "000000";
				when "000111101001011110" => data <= "000000";
				when "000111101001011111" => data <= "000000";
				when "000111101001100000" => data <= "000000";
				when "000111101001100001" => data <= "000000";
				when "000111101001100010" => data <= "000000";
				when "000111101001100011" => data <= "000000";
				when "000111101001100100" => data <= "000000";
				when "000111101001100101" => data <= "000000";
				when "000111101001100110" => data <= "000000";
				when "000111101001100111" => data <= "000000";
				when "000111101001101000" => data <= "000000";
				when "000111101001101001" => data <= "000000";
				when "000111101001101010" => data <= "000000";
				when "000111101001101011" => data <= "000000";
				when "000111101001101100" => data <= "000000";
				when "000111101001101101" => data <= "000000";
				when "000111101001101110" => data <= "000000";
				when "000111101001101111" => data <= "000000";
				when "000111101001110000" => data <= "000000";
				when "000111101001110001" => data <= "000000";
				when "000111101001110010" => data <= "000000";
				when "000111101001110011" => data <= "000000";
				when "000111101001110100" => data <= "000000";
				when "000111101001110101" => data <= "000000";
				when "000111101001110110" => data <= "000000";
				when "000111101001110111" => data <= "000000";
				when "000111101001111000" => data <= "000000";
				when "000111101001111001" => data <= "000000";
				when "000111101001111010" => data <= "000000";
				when "000111101001111011" => data <= "000000";
				when "000111101001111100" => data <= "000000";
				when "000111101001111101" => data <= "000000";
				when "000111101001111110" => data <= "000000";
				when "000111101001111111" => data <= "000000";
				when "000111101010000000" => data <= "000000";
				when "000111101010000001" => data <= "000000";
				when "000111101010000010" => data <= "000000";
				when "000111101010000011" => data <= "000000";
				when "000111101010000100" => data <= "000000";
				when "000111101010000101" => data <= "000000";
				when "000111101010000110" => data <= "000000";
				when "000111101010000111" => data <= "000000";
				when "000111101010001000" => data <= "000000";
				when "000111101010001001" => data <= "000000";
				when "000111101010001010" => data <= "000000";
				when "000111101010001011" => data <= "000000";
				when "000111101010001100" => data <= "000000";
				when "000111101010001101" => data <= "000000";
				when "000111101010001110" => data <= "000000";
				when "000111101010001111" => data <= "000000";
				when "000111101010010000" => data <= "000000";
				when "000111101010010001" => data <= "000000";
				when "000111101010010010" => data <= "000000";
				when "000111101010010011" => data <= "000000";
				when "000111101010010100" => data <= "000000";
				when "000111101010010101" => data <= "000000";
				when "000111101010010110" => data <= "000000";
				when "000111101010010111" => data <= "000000";
				when "000111101010011000" => data <= "000000";
				when "000111101010011001" => data <= "000000";
				when "000111101010011010" => data <= "000000";
				when "000111101010011011" => data <= "000000";
				when "000111101010011100" => data <= "000000";
				when "000111101010011101" => data <= "000000";
				when "000111101010011110" => data <= "000000";
				when "000111101010011111" => data <= "000000";
				when "000111110000000000" => data <= "000000";
				when "000111110000000001" => data <= "000000";
				when "000111110000000010" => data <= "000000";
				when "000111110000000011" => data <= "000000";
				when "000111110000000100" => data <= "000000";
				when "000111110000000101" => data <= "000000";
				when "000111110000000110" => data <= "000000";
				when "000111110000000111" => data <= "000000";
				when "000111110000001000" => data <= "000000";
				when "000111110000001001" => data <= "000000";
				when "000111110000001010" => data <= "000000";
				when "000111110000001011" => data <= "000000";
				when "000111110000001100" => data <= "000000";
				when "000111110000001101" => data <= "000000";
				when "000111110000001110" => data <= "000000";
				when "000111110000001111" => data <= "000000";
				when "000111110000010000" => data <= "000000";
				when "000111110000010001" => data <= "000000";
				when "000111110000010010" => data <= "000000";
				when "000111110000010011" => data <= "000000";
				when "000111110000010100" => data <= "000000";
				when "000111110000010101" => data <= "000000";
				when "000111110000010110" => data <= "000000";
				when "000111110000010111" => data <= "000000";
				when "000111110000011000" => data <= "000000";
				when "000111110000011001" => data <= "000000";
				when "000111110000011010" => data <= "000000";
				when "000111110000011011" => data <= "000000";
				when "000111110000011100" => data <= "000000";
				when "000111110000011101" => data <= "000000";
				when "000111110000011110" => data <= "000000";
				when "000111110000011111" => data <= "000000";
				when "000111110000100000" => data <= "000000";
				when "000111110000100001" => data <= "000000";
				when "000111110000100010" => data <= "000000";
				when "000111110000100011" => data <= "000000";
				when "000111110000100100" => data <= "000000";
				when "000111110000100101" => data <= "000000";
				when "000111110000100110" => data <= "000000";
				when "000111110000100111" => data <= "000000";
				when "000111110000101000" => data <= "000000";
				when "000111110000101001" => data <= "000000";
				when "000111110000101010" => data <= "000000";
				when "000111110000101011" => data <= "000000";
				when "000111110000101100" => data <= "000000";
				when "000111110000101101" => data <= "000000";
				when "000111110000101110" => data <= "000000";
				when "000111110000101111" => data <= "000000";
				when "000111110000110000" => data <= "000000";
				when "000111110000110001" => data <= "000000";
				when "000111110000110010" => data <= "000000";
				when "000111110000110011" => data <= "000000";
				when "000111110000110100" => data <= "000000";
				when "000111110000110101" => data <= "000000";
				when "000111110000110110" => data <= "000000";
				when "000111110000110111" => data <= "000000";
				when "000111110000111000" => data <= "000000";
				when "000111110000111001" => data <= "000000";
				when "000111110000111010" => data <= "000000";
				when "000111110000111011" => data <= "000000";
				when "000111110000111100" => data <= "000000";
				when "000111110000111101" => data <= "000000";
				when "000111110000111110" => data <= "000000";
				when "000111110000111111" => data <= "000000";
				when "000111110001000000" => data <= "000000";
				when "000111110001000001" => data <= "000000";
				when "000111110001000010" => data <= "000000";
				when "000111110001000011" => data <= "000000";
				when "000111110001000100" => data <= "000000";
				when "000111110001000101" => data <= "000000";
				when "000111110001000110" => data <= "000000";
				when "000111110001000111" => data <= "000000";
				when "000111110001001000" => data <= "000000";
				when "000111110001001001" => data <= "000000";
				when "000111110001001010" => data <= "000000";
				when "000111110001001011" => data <= "000000";
				when "000111110001001100" => data <= "000000";
				when "000111110001001101" => data <= "000000";
				when "000111110001001110" => data <= "000000";
				when "000111110001001111" => data <= "000000";
				when "000111110001010000" => data <= "000000";
				when "000111110001010001" => data <= "000000";
				when "000111110001010010" => data <= "000000";
				when "000111110001010011" => data <= "000000";
				when "000111110001010100" => data <= "000000";
				when "000111110001010101" => data <= "000000";
				when "000111110001010110" => data <= "000000";
				when "000111110001010111" => data <= "000000";
				when "000111110001011000" => data <= "000000";
				when "000111110001011001" => data <= "000000";
				when "000111110001011010" => data <= "000000";
				when "000111110001011011" => data <= "000000";
				when "000111110001011100" => data <= "000000";
				when "000111110001011101" => data <= "000000";
				when "000111110001011110" => data <= "000000";
				when "000111110001011111" => data <= "000000";
				when "000111110001100000" => data <= "000000";
				when "000111110001100001" => data <= "000000";
				when "000111110001100010" => data <= "000000";
				when "000111110001100011" => data <= "000000";
				when "000111110001100100" => data <= "000000";
				when "000111110001100101" => data <= "000000";
				when "000111110001100110" => data <= "000000";
				when "000111110001100111" => data <= "000000";
				when "000111110001101000" => data <= "000000";
				when "000111110001101001" => data <= "000000";
				when "000111110001101010" => data <= "000000";
				when "000111110001101011" => data <= "000000";
				when "000111110001101100" => data <= "000000";
				when "000111110001101101" => data <= "000000";
				when "000111110001101110" => data <= "000000";
				when "000111110001101111" => data <= "000000";
				when "000111110001110000" => data <= "000000";
				when "000111110001110001" => data <= "000000";
				when "000111110001110010" => data <= "000000";
				when "000111110001110011" => data <= "000000";
				when "000111110001110100" => data <= "000000";
				when "000111110001110101" => data <= "000000";
				when "000111110001110110" => data <= "000000";
				when "000111110001110111" => data <= "000000";
				when "000111110001111000" => data <= "000000";
				when "000111110001111001" => data <= "000000";
				when "000111110001111010" => data <= "000000";
				when "000111110001111011" => data <= "000000";
				when "000111110001111100" => data <= "000000";
				when "000111110001111101" => data <= "000000";
				when "000111110001111110" => data <= "000000";
				when "000111110001111111" => data <= "000000";
				when "000111110010000000" => data <= "000000";
				when "000111110010000001" => data <= "000000";
				when "000111110010000010" => data <= "000000";
				when "000111110010000011" => data <= "000000";
				when "000111110010000100" => data <= "000000";
				when "000111110010000101" => data <= "000000";
				when "000111110010000110" => data <= "000000";
				when "000111110010000111" => data <= "000000";
				when "000111110010001000" => data <= "000000";
				when "000111110010001001" => data <= "000000";
				when "000111110010001010" => data <= "000000";
				when "000111110010001011" => data <= "000000";
				when "000111110010001100" => data <= "000000";
				when "000111110010001101" => data <= "000000";
				when "000111110010001110" => data <= "000000";
				when "000111110010001111" => data <= "000000";
				when "000111110010010000" => data <= "000000";
				when "000111110010010001" => data <= "000000";
				when "000111110010010010" => data <= "000000";
				when "000111110010010011" => data <= "000000";
				when "000111110010010100" => data <= "000000";
				when "000111110010010101" => data <= "000000";
				when "000111110010010110" => data <= "000000";
				when "000111110010010111" => data <= "000000";
				when "000111110010011000" => data <= "000000";
				when "000111110010011001" => data <= "000000";
				when "000111110010011010" => data <= "000000";
				when "000111110010011011" => data <= "000000";
				when "000111110010011100" => data <= "000000";
				when "000111110010011101" => data <= "000000";
				when "000111110010011110" => data <= "000000";
				when "000111110010011111" => data <= "000000";
				when "000111111000000000" => data <= "000000";
				when "000111111000000001" => data <= "000000";
				when "000111111000000010" => data <= "000000";
				when "000111111000000011" => data <= "000000";
				when "000111111000000100" => data <= "000000";
				when "000111111000000101" => data <= "000000";
				when "000111111000000110" => data <= "000000";
				when "000111111000000111" => data <= "000000";
				when "000111111000001000" => data <= "000000";
				when "000111111000001001" => data <= "000000";
				when "000111111000001010" => data <= "000000";
				when "000111111000001011" => data <= "000000";
				when "000111111000001100" => data <= "000000";
				when "000111111000001101" => data <= "000000";
				when "000111111000001110" => data <= "000000";
				when "000111111000001111" => data <= "000000";
				when "000111111000010000" => data <= "000000";
				when "000111111000010001" => data <= "000000";
				when "000111111000010010" => data <= "000000";
				when "000111111000010011" => data <= "000000";
				when "000111111000010100" => data <= "000000";
				when "000111111000010101" => data <= "000000";
				when "000111111000010110" => data <= "000000";
				when "000111111000010111" => data <= "000000";
				when "000111111000011000" => data <= "000000";
				when "000111111000011001" => data <= "000000";
				when "000111111000011010" => data <= "000000";
				when "000111111000011011" => data <= "000000";
				when "000111111000011100" => data <= "000000";
				when "000111111000011101" => data <= "000000";
				when "000111111000011110" => data <= "000000";
				when "000111111000011111" => data <= "000000";
				when "000111111000100000" => data <= "000000";
				when "000111111000100001" => data <= "000000";
				when "000111111000100010" => data <= "000000";
				when "000111111000100011" => data <= "000000";
				when "000111111000100100" => data <= "000000";
				when "000111111000100101" => data <= "000000";
				when "000111111000100110" => data <= "000000";
				when "000111111000100111" => data <= "000000";
				when "000111111000101000" => data <= "000000";
				when "000111111000101001" => data <= "000000";
				when "000111111000101010" => data <= "000000";
				when "000111111000101011" => data <= "000000";
				when "000111111000101100" => data <= "000000";
				when "000111111000101101" => data <= "000000";
				when "000111111000101110" => data <= "000000";
				when "000111111000101111" => data <= "000000";
				when "000111111000110000" => data <= "000000";
				when "000111111000110001" => data <= "000000";
				when "000111111000110010" => data <= "000000";
				when "000111111000110011" => data <= "000000";
				when "000111111000110100" => data <= "000000";
				when "000111111000110101" => data <= "000000";
				when "000111111000110110" => data <= "000000";
				when "000111111000110111" => data <= "000000";
				when "000111111000111000" => data <= "000000";
				when "000111111000111001" => data <= "000000";
				when "000111111000111010" => data <= "000000";
				when "000111111000111011" => data <= "000000";
				when "000111111000111100" => data <= "000000";
				when "000111111000111101" => data <= "000000";
				when "000111111000111110" => data <= "000000";
				when "000111111000111111" => data <= "000000";
				when "000111111001000000" => data <= "000000";
				when "000111111001000001" => data <= "000000";
				when "000111111001000010" => data <= "000000";
				when "000111111001000011" => data <= "000000";
				when "000111111001000100" => data <= "000000";
				when "000111111001000101" => data <= "000000";
				when "000111111001000110" => data <= "000000";
				when "000111111001000111" => data <= "000000";
				when "000111111001001000" => data <= "000000";
				when "000111111001001001" => data <= "000000";
				when "000111111001001010" => data <= "000000";
				when "000111111001001011" => data <= "000000";
				when "000111111001001100" => data <= "000000";
				when "000111111001001101" => data <= "000000";
				when "000111111001001110" => data <= "000000";
				when "000111111001001111" => data <= "000000";
				when "000111111001010000" => data <= "000000";
				when "000111111001010001" => data <= "000000";
				when "000111111001010010" => data <= "000000";
				when "000111111001010011" => data <= "000000";
				when "000111111001010100" => data <= "000000";
				when "000111111001010101" => data <= "000000";
				when "000111111001010110" => data <= "000000";
				when "000111111001010111" => data <= "000000";
				when "000111111001011000" => data <= "000000";
				when "000111111001011001" => data <= "000000";
				when "000111111001011010" => data <= "000000";
				when "000111111001011011" => data <= "000000";
				when "000111111001011100" => data <= "000000";
				when "000111111001011101" => data <= "000000";
				when "000111111001011110" => data <= "000000";
				when "000111111001011111" => data <= "000000";
				when "000111111001100000" => data <= "000000";
				when "000111111001100001" => data <= "000000";
				when "000111111001100010" => data <= "000000";
				when "000111111001100011" => data <= "000000";
				when "000111111001100100" => data <= "000000";
				when "000111111001100101" => data <= "000000";
				when "000111111001100110" => data <= "000000";
				when "000111111001100111" => data <= "000000";
				when "000111111001101000" => data <= "000000";
				when "000111111001101001" => data <= "000000";
				when "000111111001101010" => data <= "000000";
				when "000111111001101011" => data <= "000000";
				when "000111111001101100" => data <= "000000";
				when "000111111001101101" => data <= "000000";
				when "000111111001101110" => data <= "000000";
				when "000111111001101111" => data <= "000000";
				when "000111111001110000" => data <= "000000";
				when "000111111001110001" => data <= "000000";
				when "000111111001110010" => data <= "000000";
				when "000111111001110011" => data <= "000000";
				when "000111111001110100" => data <= "000000";
				when "000111111001110101" => data <= "000000";
				when "000111111001110110" => data <= "000000";
				when "000111111001110111" => data <= "000000";
				when "000111111001111000" => data <= "000000";
				when "000111111001111001" => data <= "000000";
				when "000111111001111010" => data <= "000000";
				when "000111111001111011" => data <= "000000";
				when "000111111001111100" => data <= "000000";
				when "000111111001111101" => data <= "000000";
				when "000111111001111110" => data <= "000000";
				when "000111111001111111" => data <= "000000";
				when "000111111010000000" => data <= "000000";
				when "000111111010000001" => data <= "000000";
				when "000111111010000010" => data <= "000000";
				when "000111111010000011" => data <= "000000";
				when "000111111010000100" => data <= "000000";
				when "000111111010000101" => data <= "000000";
				when "000111111010000110" => data <= "000000";
				when "000111111010000111" => data <= "000000";
				when "000111111010001000" => data <= "000000";
				when "000111111010001001" => data <= "000000";
				when "000111111010001010" => data <= "000000";
				when "000111111010001011" => data <= "000000";
				when "000111111010001100" => data <= "000000";
				when "000111111010001101" => data <= "000000";
				when "000111111010001110" => data <= "000000";
				when "000111111010001111" => data <= "000000";
				when "000111111010010000" => data <= "000000";
				when "000111111010010001" => data <= "000000";
				when "000111111010010010" => data <= "000000";
				when "000111111010010011" => data <= "000000";
				when "000111111010010100" => data <= "000000";
				when "000111111010010101" => data <= "000000";
				when "000111111010010110" => data <= "000000";
				when "000111111010010111" => data <= "000000";
				when "000111111010011000" => data <= "000000";
				when "000111111010011001" => data <= "000000";
				when "000111111010011010" => data <= "000000";
				when "000111111010011011" => data <= "000000";
				when "000111111010011100" => data <= "000000";
				when "000111111010011101" => data <= "000000";
				when "000111111010011110" => data <= "000000";
				when "000111111010011111" => data <= "000000";
				when "001000000000000000" => data <= "000000";
				when "001000000000000001" => data <= "000000";
				when "001000000000000010" => data <= "000000";
				when "001000000000000011" => data <= "000000";
				when "001000000000000100" => data <= "000000";
				when "001000000000000101" => data <= "000000";
				when "001000000000000110" => data <= "000000";
				when "001000000000000111" => data <= "000000";
				when "001000000000001000" => data <= "000000";
				when "001000000000001001" => data <= "000000";
				when "001000000000001010" => data <= "000000";
				when "001000000000001011" => data <= "000000";
				when "001000000000001100" => data <= "000000";
				when "001000000000001101" => data <= "000000";
				when "001000000000001110" => data <= "000000";
				when "001000000000001111" => data <= "000000";
				when "001000000000010000" => data <= "000000";
				when "001000000000010001" => data <= "000000";
				when "001000000000010010" => data <= "000000";
				when "001000000000010011" => data <= "000000";
				when "001000000000010100" => data <= "000000";
				when "001000000000010101" => data <= "000000";
				when "001000000000010110" => data <= "000000";
				when "001000000000010111" => data <= "000000";
				when "001000000000011000" => data <= "000000";
				when "001000000000011001" => data <= "000000";
				when "001000000000011010" => data <= "000000";
				when "001000000000011011" => data <= "000000";
				when "001000000000011100" => data <= "000000";
				when "001000000000011101" => data <= "000000";
				when "001000000000011110" => data <= "000000";
				when "001000000000011111" => data <= "000000";
				when "001000000000100000" => data <= "000000";
				when "001000000000100001" => data <= "000000";
				when "001000000000100010" => data <= "000000";
				when "001000000000100011" => data <= "000000";
				when "001000000000100100" => data <= "000000";
				when "001000000000100101" => data <= "000000";
				when "001000000000100110" => data <= "000000";
				when "001000000000100111" => data <= "000000";
				when "001000000000101000" => data <= "000000";
				when "001000000000101001" => data <= "000000";
				when "001000000000101010" => data <= "000000";
				when "001000000000101011" => data <= "000000";
				when "001000000000101100" => data <= "000000";
				when "001000000000101101" => data <= "000000";
				when "001000000000101110" => data <= "000000";
				when "001000000000101111" => data <= "000000";
				when "001000000000110000" => data <= "000000";
				when "001000000000110001" => data <= "000000";
				when "001000000000110010" => data <= "000000";
				when "001000000000110011" => data <= "000000";
				when "001000000000110100" => data <= "000000";
				when "001000000000110101" => data <= "000000";
				when "001000000000110110" => data <= "000000";
				when "001000000000110111" => data <= "000000";
				when "001000000000111000" => data <= "000000";
				when "001000000000111001" => data <= "000000";
				when "001000000000111010" => data <= "000000";
				when "001000000000111011" => data <= "000000";
				when "001000000000111100" => data <= "000000";
				when "001000000000111101" => data <= "000000";
				when "001000000000111110" => data <= "000000";
				when "001000000000111111" => data <= "000000";
				when "001000000001000000" => data <= "000000";
				when "001000000001000001" => data <= "000000";
				when "001000000001000010" => data <= "000000";
				when "001000000001000011" => data <= "000000";
				when "001000000001000100" => data <= "000000";
				when "001000000001000101" => data <= "000000";
				when "001000000001000110" => data <= "000000";
				when "001000000001000111" => data <= "000000";
				when "001000000001001000" => data <= "000000";
				when "001000000001001001" => data <= "000000";
				when "001000000001001010" => data <= "000000";
				when "001000000001001011" => data <= "000000";
				when "001000000001001100" => data <= "000000";
				when "001000000001001101" => data <= "000000";
				when "001000000001001110" => data <= "000000";
				when "001000000001001111" => data <= "000000";
				when "001000000001010000" => data <= "000000";
				when "001000000001010001" => data <= "000000";
				when "001000000001010010" => data <= "000000";
				when "001000000001010011" => data <= "000000";
				when "001000000001010100" => data <= "000000";
				when "001000000001010101" => data <= "000000";
				when "001000000001010110" => data <= "000000";
				when "001000000001010111" => data <= "000000";
				when "001000000001011000" => data <= "000000";
				when "001000000001011001" => data <= "000000";
				when "001000000001011010" => data <= "000000";
				when "001000000001011011" => data <= "000000";
				when "001000000001011100" => data <= "000000";
				when "001000000001011101" => data <= "000000";
				when "001000000001011110" => data <= "000000";
				when "001000000001011111" => data <= "000000";
				when "001000000001100000" => data <= "000000";
				when "001000000001100001" => data <= "000000";
				when "001000000001100010" => data <= "000000";
				when "001000000001100011" => data <= "000000";
				when "001000000001100100" => data <= "000000";
				when "001000000001100101" => data <= "000000";
				when "001000000001100110" => data <= "000000";
				when "001000000001100111" => data <= "000000";
				when "001000000001101000" => data <= "000000";
				when "001000000001101001" => data <= "000000";
				when "001000000001101010" => data <= "000000";
				when "001000000001101011" => data <= "000000";
				when "001000000001101100" => data <= "000000";
				when "001000000001101101" => data <= "000000";
				when "001000000001101110" => data <= "000000";
				when "001000000001101111" => data <= "000000";
				when "001000000001110000" => data <= "000000";
				when "001000000001110001" => data <= "000000";
				when "001000000001110010" => data <= "000000";
				when "001000000001110011" => data <= "000000";
				when "001000000001110100" => data <= "000000";
				when "001000000001110101" => data <= "000000";
				when "001000000001110110" => data <= "000000";
				when "001000000001110111" => data <= "000000";
				when "001000000001111000" => data <= "000000";
				when "001000000001111001" => data <= "000000";
				when "001000000001111010" => data <= "000000";
				when "001000000001111011" => data <= "000000";
				when "001000000001111100" => data <= "000000";
				when "001000000001111101" => data <= "000000";
				when "001000000001111110" => data <= "000000";
				when "001000000001111111" => data <= "000000";
				when "001000000010000000" => data <= "000000";
				when "001000000010000001" => data <= "000000";
				when "001000000010000010" => data <= "000000";
				when "001000000010000011" => data <= "000000";
				when "001000000010000100" => data <= "000000";
				when "001000000010000101" => data <= "000000";
				when "001000000010000110" => data <= "000000";
				when "001000000010000111" => data <= "000000";
				when "001000000010001000" => data <= "000000";
				when "001000000010001001" => data <= "000000";
				when "001000000010001010" => data <= "000000";
				when "001000000010001011" => data <= "000000";
				when "001000000010001100" => data <= "000000";
				when "001000000010001101" => data <= "000000";
				when "001000000010001110" => data <= "000000";
				when "001000000010001111" => data <= "000000";
				when "001000000010010000" => data <= "000000";
				when "001000000010010001" => data <= "000000";
				when "001000000010010010" => data <= "000000";
				when "001000000010010011" => data <= "000000";
				when "001000000010010100" => data <= "000000";
				when "001000000010010101" => data <= "000000";
				when "001000000010010110" => data <= "000000";
				when "001000000010010111" => data <= "000000";
				when "001000000010011000" => data <= "000000";
				when "001000000010011001" => data <= "000000";
				when "001000000010011010" => data <= "000000";
				when "001000000010011011" => data <= "000000";
				when "001000000010011100" => data <= "000000";
				when "001000000010011101" => data <= "000000";
				when "001000000010011110" => data <= "000000";
				when "001000000010011111" => data <= "000000";
				when "001000001000000000" => data <= "000000";
				when "001000001000000001" => data <= "000000";
				when "001000001000000010" => data <= "000000";
				when "001000001000000011" => data <= "000000";
				when "001000001000000100" => data <= "000000";
				when "001000001000000101" => data <= "000000";
				when "001000001000000110" => data <= "000000";
				when "001000001000000111" => data <= "000000";
				when "001000001000001000" => data <= "000000";
				when "001000001000001001" => data <= "000000";
				when "001000001000001010" => data <= "000000";
				when "001000001000001011" => data <= "000000";
				when "001000001000001100" => data <= "000000";
				when "001000001000001101" => data <= "000000";
				when "001000001000001110" => data <= "000000";
				when "001000001000001111" => data <= "000000";
				when "001000001000010000" => data <= "000000";
				when "001000001000010001" => data <= "000000";
				when "001000001000010010" => data <= "000000";
				when "001000001000010011" => data <= "000000";
				when "001000001000010100" => data <= "000000";
				when "001000001000010101" => data <= "000000";
				when "001000001000010110" => data <= "000000";
				when "001000001000010111" => data <= "000000";
				when "001000001000011000" => data <= "000000";
				when "001000001000011001" => data <= "000000";
				when "001000001000011010" => data <= "000000";
				when "001000001000011011" => data <= "000000";
				when "001000001000011100" => data <= "000000";
				when "001000001000011101" => data <= "000000";
				when "001000001000011110" => data <= "000000";
				when "001000001000011111" => data <= "000000";
				when "001000001000100000" => data <= "000000";
				when "001000001000100001" => data <= "000000";
				when "001000001000100010" => data <= "000000";
				when "001000001000100011" => data <= "000000";
				when "001000001000100100" => data <= "000000";
				when "001000001000100101" => data <= "000000";
				when "001000001000100110" => data <= "000000";
				when "001000001000100111" => data <= "000000";
				when "001000001000101000" => data <= "000000";
				when "001000001000101001" => data <= "000000";
				when "001000001000101010" => data <= "000000";
				when "001000001000101011" => data <= "000000";
				when "001000001000101100" => data <= "000000";
				when "001000001000101101" => data <= "000000";
				when "001000001000101110" => data <= "000000";
				when "001000001000101111" => data <= "000000";
				when "001000001000110000" => data <= "000000";
				when "001000001000110001" => data <= "000000";
				when "001000001000110010" => data <= "000000";
				when "001000001000110011" => data <= "000000";
				when "001000001000110100" => data <= "000000";
				when "001000001000110101" => data <= "000000";
				when "001000001000110110" => data <= "000000";
				when "001000001000110111" => data <= "000000";
				when "001000001000111000" => data <= "000000";
				when "001000001000111001" => data <= "000000";
				when "001000001000111010" => data <= "000000";
				when "001000001000111011" => data <= "000000";
				when "001000001000111100" => data <= "000000";
				when "001000001000111101" => data <= "000000";
				when "001000001000111110" => data <= "000000";
				when "001000001000111111" => data <= "000000";
				when "001000001001000000" => data <= "000000";
				when "001000001001000001" => data <= "000000";
				when "001000001001000010" => data <= "000000";
				when "001000001001000011" => data <= "000000";
				when "001000001001000100" => data <= "000000";
				when "001000001001000101" => data <= "000000";
				when "001000001001000110" => data <= "000000";
				when "001000001001000111" => data <= "000000";
				when "001000001001001000" => data <= "000000";
				when "001000001001001001" => data <= "000000";
				when "001000001001001010" => data <= "000000";
				when "001000001001001011" => data <= "000000";
				when "001000001001001100" => data <= "000000";
				when "001000001001001101" => data <= "000000";
				when "001000001001001110" => data <= "000000";
				when "001000001001001111" => data <= "000000";
				when "001000001001010000" => data <= "000000";
				when "001000001001010001" => data <= "000000";
				when "001000001001010010" => data <= "000000";
				when "001000001001010011" => data <= "000000";
				when "001000001001010100" => data <= "000000";
				when "001000001001010101" => data <= "000000";
				when "001000001001010110" => data <= "000000";
				when "001000001001010111" => data <= "000000";
				when "001000001001011000" => data <= "000000";
				when "001000001001011001" => data <= "000000";
				when "001000001001011010" => data <= "000000";
				when "001000001001011011" => data <= "000000";
				when "001000001001011100" => data <= "000000";
				when "001000001001011101" => data <= "000000";
				when "001000001001011110" => data <= "000000";
				when "001000001001011111" => data <= "000000";
				when "001000001001100000" => data <= "000000";
				when "001000001001100001" => data <= "000000";
				when "001000001001100010" => data <= "000000";
				when "001000001001100011" => data <= "000000";
				when "001000001001100100" => data <= "000000";
				when "001000001001100101" => data <= "000000";
				when "001000001001100110" => data <= "000000";
				when "001000001001100111" => data <= "000000";
				when "001000001001101000" => data <= "000000";
				when "001000001001101001" => data <= "000000";
				when "001000001001101010" => data <= "000000";
				when "001000001001101011" => data <= "000000";
				when "001000001001101100" => data <= "000000";
				when "001000001001101101" => data <= "000000";
				when "001000001001101110" => data <= "000000";
				when "001000001001101111" => data <= "000000";
				when "001000001001110000" => data <= "000000";
				when "001000001001110001" => data <= "000000";
				when "001000001001110010" => data <= "000000";
				when "001000001001110011" => data <= "000000";
				when "001000001001110100" => data <= "000000";
				when "001000001001110101" => data <= "000000";
				when "001000001001110110" => data <= "000000";
				when "001000001001110111" => data <= "000000";
				when "001000001001111000" => data <= "000000";
				when "001000001001111001" => data <= "000000";
				when "001000001001111010" => data <= "000000";
				when "001000001001111011" => data <= "000000";
				when "001000001001111100" => data <= "000000";
				when "001000001001111101" => data <= "000000";
				when "001000001001111110" => data <= "000000";
				when "001000001001111111" => data <= "000000";
				when "001000001010000000" => data <= "000000";
				when "001000001010000001" => data <= "000000";
				when "001000001010000010" => data <= "000000";
				when "001000001010000011" => data <= "000000";
				when "001000001010000100" => data <= "000000";
				when "001000001010000101" => data <= "000000";
				when "001000001010000110" => data <= "000000";
				when "001000001010000111" => data <= "000000";
				when "001000001010001000" => data <= "000000";
				when "001000001010001001" => data <= "000000";
				when "001000001010001010" => data <= "000000";
				when "001000001010001011" => data <= "000000";
				when "001000001010001100" => data <= "000000";
				when "001000001010001101" => data <= "000000";
				when "001000001010001110" => data <= "000000";
				when "001000001010001111" => data <= "000000";
				when "001000001010010000" => data <= "000000";
				when "001000001010010001" => data <= "000000";
				when "001000001010010010" => data <= "000000";
				when "001000001010010011" => data <= "000000";
				when "001000001010010100" => data <= "000000";
				when "001000001010010101" => data <= "000000";
				when "001000001010010110" => data <= "000000";
				when "001000001010010111" => data <= "000000";
				when "001000001010011000" => data <= "000000";
				when "001000001010011001" => data <= "000000";
				when "001000001010011010" => data <= "000000";
				when "001000001010011011" => data <= "000000";
				when "001000001010011100" => data <= "000000";
				when "001000001010011101" => data <= "000000";
				when "001000001010011110" => data <= "000000";
				when "001000001010011111" => data <= "000000";
				when "001000010000000000" => data <= "000000";
				when "001000010000000001" => data <= "000000";
				when "001000010000000010" => data <= "000000";
				when "001000010000000011" => data <= "000000";
				when "001000010000000100" => data <= "000000";
				when "001000010000000101" => data <= "000000";
				when "001000010000000110" => data <= "000000";
				when "001000010000000111" => data <= "000000";
				when "001000010000001000" => data <= "000000";
				when "001000010000001001" => data <= "000000";
				when "001000010000001010" => data <= "000000";
				when "001000010000001011" => data <= "000000";
				when "001000010000001100" => data <= "000000";
				when "001000010000001101" => data <= "000000";
				when "001000010000001110" => data <= "000000";
				when "001000010000001111" => data <= "000000";
				when "001000010000010000" => data <= "000000";
				when "001000010000010001" => data <= "000000";
				when "001000010000010010" => data <= "000000";
				when "001000010000010011" => data <= "000000";
				when "001000010000010100" => data <= "000000";
				when "001000010000010101" => data <= "000000";
				when "001000010000010110" => data <= "000000";
				when "001000010000010111" => data <= "000000";
				when "001000010000011000" => data <= "000000";
				when "001000010000011001" => data <= "000000";
				when "001000010000011010" => data <= "000000";
				when "001000010000011011" => data <= "000000";
				when "001000010000011100" => data <= "000000";
				when "001000010000011101" => data <= "000000";
				when "001000010000011110" => data <= "000000";
				when "001000010000011111" => data <= "000000";
				when "001000010000100000" => data <= "000000";
				when "001000010000100001" => data <= "000000";
				when "001000010000100010" => data <= "000000";
				when "001000010000100011" => data <= "000000";
				when "001000010000100100" => data <= "000000";
				when "001000010000100101" => data <= "000000";
				when "001000010000100110" => data <= "000000";
				when "001000010000100111" => data <= "000000";
				when "001000010000101000" => data <= "000000";
				when "001000010000101001" => data <= "000000";
				when "001000010000101010" => data <= "000000";
				when "001000010000101011" => data <= "000000";
				when "001000010000101100" => data <= "000000";
				when "001000010000101101" => data <= "000000";
				when "001000010000101110" => data <= "000000";
				when "001000010000101111" => data <= "000000";
				when "001000010000110000" => data <= "000000";
				when "001000010000110001" => data <= "000000";
				when "001000010000110010" => data <= "000000";
				when "001000010000110011" => data <= "000000";
				when "001000010000110100" => data <= "000000";
				when "001000010000110101" => data <= "000000";
				when "001000010000110110" => data <= "000000";
				when "001000010000110111" => data <= "000000";
				when "001000010000111000" => data <= "000000";
				when "001000010000111001" => data <= "000000";
				when "001000010000111010" => data <= "000000";
				when "001000010000111011" => data <= "000000";
				when "001000010000111100" => data <= "000000";
				when "001000010000111101" => data <= "000000";
				when "001000010000111110" => data <= "000000";
				when "001000010000111111" => data <= "000000";
				when "001000010001000000" => data <= "000000";
				when "001000010001000001" => data <= "000000";
				when "001000010001000010" => data <= "000000";
				when "001000010001000011" => data <= "000000";
				when "001000010001000100" => data <= "000000";
				when "001000010001000101" => data <= "000000";
				when "001000010001000110" => data <= "000000";
				when "001000010001000111" => data <= "000000";
				when "001000010001001000" => data <= "000000";
				when "001000010001001001" => data <= "000000";
				when "001000010001001010" => data <= "000000";
				when "001000010001001011" => data <= "000000";
				when "001000010001001100" => data <= "000000";
				when "001000010001001101" => data <= "000000";
				when "001000010001001110" => data <= "000000";
				when "001000010001001111" => data <= "000000";
				when "001000010001010000" => data <= "000000";
				when "001000010001010001" => data <= "000000";
				when "001000010001010010" => data <= "000000";
				when "001000010001010011" => data <= "000000";
				when "001000010001010100" => data <= "000000";
				when "001000010001010101" => data <= "000000";
				when "001000010001010110" => data <= "000000";
				when "001000010001010111" => data <= "000000";
				when "001000010001011000" => data <= "000000";
				when "001000010001011001" => data <= "000000";
				when "001000010001011010" => data <= "000000";
				when "001000010001011011" => data <= "000000";
				when "001000010001011100" => data <= "000000";
				when "001000010001011101" => data <= "000000";
				when "001000010001011110" => data <= "000000";
				when "001000010001011111" => data <= "000000";
				when "001000010001100000" => data <= "000000";
				when "001000010001100001" => data <= "000000";
				when "001000010001100010" => data <= "000000";
				when "001000010001100011" => data <= "000000";
				when "001000010001100100" => data <= "000000";
				when "001000010001100101" => data <= "000000";
				when "001000010001100110" => data <= "000000";
				when "001000010001100111" => data <= "000000";
				when "001000010001101000" => data <= "000000";
				when "001000010001101001" => data <= "000000";
				when "001000010001101010" => data <= "000000";
				when "001000010001101011" => data <= "000000";
				when "001000010001101100" => data <= "000000";
				when "001000010001101101" => data <= "000000";
				when "001000010001101110" => data <= "000000";
				when "001000010001101111" => data <= "000000";
				when "001000010001110000" => data <= "000000";
				when "001000010001110001" => data <= "000000";
				when "001000010001110010" => data <= "000000";
				when "001000010001110011" => data <= "000000";
				when "001000010001110100" => data <= "000000";
				when "001000010001110101" => data <= "000000";
				when "001000010001110110" => data <= "000000";
				when "001000010001110111" => data <= "000000";
				when "001000010001111000" => data <= "000000";
				when "001000010001111001" => data <= "000000";
				when "001000010001111010" => data <= "000000";
				when "001000010001111011" => data <= "000000";
				when "001000010001111100" => data <= "000000";
				when "001000010001111101" => data <= "000000";
				when "001000010001111110" => data <= "000000";
				when "001000010001111111" => data <= "000000";
				when "001000010010000000" => data <= "000000";
				when "001000010010000001" => data <= "000000";
				when "001000010010000010" => data <= "000000";
				when "001000010010000011" => data <= "000000";
				when "001000010010000100" => data <= "000000";
				when "001000010010000101" => data <= "000000";
				when "001000010010000110" => data <= "000000";
				when "001000010010000111" => data <= "000000";
				when "001000010010001000" => data <= "000000";
				when "001000010010001001" => data <= "000000";
				when "001000010010001010" => data <= "000000";
				when "001000010010001011" => data <= "000000";
				when "001000010010001100" => data <= "000000";
				when "001000010010001101" => data <= "000000";
				when "001000010010001110" => data <= "000000";
				when "001000010010001111" => data <= "000000";
				when "001000010010010000" => data <= "000000";
				when "001000010010010001" => data <= "000000";
				when "001000010010010010" => data <= "000000";
				when "001000010010010011" => data <= "000000";
				when "001000010010010100" => data <= "000000";
				when "001000010010010101" => data <= "000000";
				when "001000010010010110" => data <= "000000";
				when "001000010010010111" => data <= "000000";
				when "001000010010011000" => data <= "000000";
				when "001000010010011001" => data <= "000000";
				when "001000010010011010" => data <= "000000";
				when "001000010010011011" => data <= "000000";
				when "001000010010011100" => data <= "000000";
				when "001000010010011101" => data <= "000000";
				when "001000010010011110" => data <= "000000";
				when "001000010010011111" => data <= "000000";
				when "001000011000000000" => data <= "000000";
				when "001000011000000001" => data <= "000000";
				when "001000011000000010" => data <= "000000";
				when "001000011000000011" => data <= "000000";
				when "001000011000000100" => data <= "000000";
				when "001000011000000101" => data <= "000000";
				when "001000011000000110" => data <= "000000";
				when "001000011000000111" => data <= "000000";
				when "001000011000001000" => data <= "000000";
				when "001000011000001001" => data <= "000000";
				when "001000011000001010" => data <= "000000";
				when "001000011000001011" => data <= "000000";
				when "001000011000001100" => data <= "000000";
				when "001000011000001101" => data <= "000000";
				when "001000011000001110" => data <= "000000";
				when "001000011000001111" => data <= "000000";
				when "001000011000010000" => data <= "000000";
				when "001000011000010001" => data <= "000000";
				when "001000011000010010" => data <= "000000";
				when "001000011000010011" => data <= "000000";
				when "001000011000010100" => data <= "000000";
				when "001000011000010101" => data <= "000000";
				when "001000011000010110" => data <= "000000";
				when "001000011000010111" => data <= "000000";
				when "001000011000011000" => data <= "000000";
				when "001000011000011001" => data <= "000000";
				when "001000011000011010" => data <= "000000";
				when "001000011000011011" => data <= "000000";
				when "001000011000011100" => data <= "000000";
				when "001000011000011101" => data <= "000000";
				when "001000011000011110" => data <= "000000";
				when "001000011000011111" => data <= "000000";
				when "001000011000100000" => data <= "000000";
				when "001000011000100001" => data <= "000000";
				when "001000011000100010" => data <= "000000";
				when "001000011000100011" => data <= "000000";
				when "001000011000100100" => data <= "000000";
				when "001000011000100101" => data <= "000000";
				when "001000011000100110" => data <= "000000";
				when "001000011000100111" => data <= "000000";
				when "001000011000101000" => data <= "000000";
				when "001000011000101001" => data <= "000000";
				when "001000011000101010" => data <= "000000";
				when "001000011000101011" => data <= "000000";
				when "001000011000101100" => data <= "000000";
				when "001000011000101101" => data <= "000000";
				when "001000011000101110" => data <= "000000";
				when "001000011000101111" => data <= "000000";
				when "001000011000110000" => data <= "000000";
				when "001000011000110001" => data <= "000000";
				when "001000011000110010" => data <= "000000";
				when "001000011000110011" => data <= "000000";
				when "001000011000110100" => data <= "000000";
				when "001000011000110101" => data <= "000000";
				when "001000011000110110" => data <= "000000";
				when "001000011000110111" => data <= "000000";
				when "001000011000111000" => data <= "000000";
				when "001000011000111001" => data <= "000000";
				when "001000011000111010" => data <= "000000";
				when "001000011000111011" => data <= "000000";
				when "001000011000111100" => data <= "000000";
				when "001000011000111101" => data <= "000000";
				when "001000011000111110" => data <= "000000";
				when "001000011000111111" => data <= "000000";
				when "001000011001000000" => data <= "000000";
				when "001000011001000001" => data <= "000000";
				when "001000011001000010" => data <= "000000";
				when "001000011001000011" => data <= "000000";
				when "001000011001000100" => data <= "000000";
				when "001000011001000101" => data <= "000000";
				when "001000011001000110" => data <= "000000";
				when "001000011001000111" => data <= "000000";
				when "001000011001001000" => data <= "000000";
				when "001000011001001001" => data <= "000000";
				when "001000011001001010" => data <= "000000";
				when "001000011001001011" => data <= "000000";
				when "001000011001001100" => data <= "000000";
				when "001000011001001101" => data <= "000000";
				when "001000011001001110" => data <= "000000";
				when "001000011001001111" => data <= "000000";
				when "001000011001010000" => data <= "000000";
				when "001000011001010001" => data <= "000000";
				when "001000011001010010" => data <= "000000";
				when "001000011001010011" => data <= "000000";
				when "001000011001010100" => data <= "000000";
				when "001000011001010101" => data <= "000000";
				when "001000011001010110" => data <= "000000";
				when "001000011001010111" => data <= "000000";
				when "001000011001011000" => data <= "000000";
				when "001000011001011001" => data <= "000000";
				when "001000011001011010" => data <= "000000";
				when "001000011001011011" => data <= "000000";
				when "001000011001011100" => data <= "000000";
				when "001000011001011101" => data <= "000000";
				when "001000011001011110" => data <= "000000";
				when "001000011001011111" => data <= "000000";
				when "001000011001100000" => data <= "000000";
				when "001000011001100001" => data <= "000000";
				when "001000011001100010" => data <= "000000";
				when "001000011001100011" => data <= "000000";
				when "001000011001100100" => data <= "000000";
				when "001000011001100101" => data <= "000000";
				when "001000011001100110" => data <= "000000";
				when "001000011001100111" => data <= "000000";
				when "001000011001101000" => data <= "000000";
				when "001000011001101001" => data <= "000000";
				when "001000011001101010" => data <= "000000";
				when "001000011001101011" => data <= "000000";
				when "001000011001101100" => data <= "000000";
				when "001000011001101101" => data <= "000000";
				when "001000011001101110" => data <= "000000";
				when "001000011001101111" => data <= "000000";
				when "001000011001110000" => data <= "000000";
				when "001000011001110001" => data <= "000000";
				when "001000011001110010" => data <= "000000";
				when "001000011001110011" => data <= "000000";
				when "001000011001110100" => data <= "000000";
				when "001000011001110101" => data <= "000000";
				when "001000011001110110" => data <= "000000";
				when "001000011001110111" => data <= "000000";
				when "001000011001111000" => data <= "000000";
				when "001000011001111001" => data <= "000000";
				when "001000011001111010" => data <= "000000";
				when "001000011001111011" => data <= "000000";
				when "001000011001111100" => data <= "000000";
				when "001000011001111101" => data <= "000000";
				when "001000011001111110" => data <= "000000";
				when "001000011001111111" => data <= "000000";
				when "001000011010000000" => data <= "000000";
				when "001000011010000001" => data <= "000000";
				when "001000011010000010" => data <= "000000";
				when "001000011010000011" => data <= "000000";
				when "001000011010000100" => data <= "000000";
				when "001000011010000101" => data <= "000000";
				when "001000011010000110" => data <= "000000";
				when "001000011010000111" => data <= "000000";
				when "001000011010001000" => data <= "000000";
				when "001000011010001001" => data <= "000000";
				when "001000011010001010" => data <= "000000";
				when "001000011010001011" => data <= "000000";
				when "001000011010001100" => data <= "000000";
				when "001000011010001101" => data <= "000000";
				when "001000011010001110" => data <= "000000";
				when "001000011010001111" => data <= "000000";
				when "001000011010010000" => data <= "000000";
				when "001000011010010001" => data <= "000000";
				when "001000011010010010" => data <= "000000";
				when "001000011010010011" => data <= "000000";
				when "001000011010010100" => data <= "000000";
				when "001000011010010101" => data <= "000000";
				when "001000011010010110" => data <= "000000";
				when "001000011010010111" => data <= "000000";
				when "001000011010011000" => data <= "000000";
				when "001000011010011001" => data <= "000000";
				when "001000011010011010" => data <= "000000";
				when "001000011010011011" => data <= "000000";
				when "001000011010011100" => data <= "000000";
				when "001000011010011101" => data <= "000000";
				when "001000011010011110" => data <= "000000";
				when "001000011010011111" => data <= "000000";
				when "001000100000000000" => data <= "000000";
				when "001000100000000001" => data <= "000000";
				when "001000100000000010" => data <= "000000";
				when "001000100000000011" => data <= "000000";
				when "001000100000000100" => data <= "000000";
				when "001000100000000101" => data <= "000000";
				when "001000100000000110" => data <= "000000";
				when "001000100000000111" => data <= "000000";
				when "001000100000001000" => data <= "000000";
				when "001000100000001001" => data <= "000000";
				when "001000100000001010" => data <= "000000";
				when "001000100000001011" => data <= "000000";
				when "001000100000001100" => data <= "000000";
				when "001000100000001101" => data <= "000000";
				when "001000100000001110" => data <= "000000";
				when "001000100000001111" => data <= "000000";
				when "001000100000010000" => data <= "000000";
				when "001000100000010001" => data <= "000000";
				when "001000100000010010" => data <= "000000";
				when "001000100000010011" => data <= "000000";
				when "001000100000010100" => data <= "000000";
				when "001000100000010101" => data <= "000000";
				when "001000100000010110" => data <= "000000";
				when "001000100000010111" => data <= "000000";
				when "001000100000011000" => data <= "000000";
				when "001000100000011001" => data <= "000000";
				when "001000100000011010" => data <= "000000";
				when "001000100000011011" => data <= "000000";
				when "001000100000011100" => data <= "000000";
				when "001000100000011101" => data <= "000000";
				when "001000100000011110" => data <= "000000";
				when "001000100000011111" => data <= "000000";
				when "001000100000100000" => data <= "000000";
				when "001000100000100001" => data <= "000000";
				when "001000100000100010" => data <= "000000";
				when "001000100000100011" => data <= "000000";
				when "001000100000100100" => data <= "000000";
				when "001000100000100101" => data <= "000000";
				when "001000100000100110" => data <= "000000";
				when "001000100000100111" => data <= "000000";
				when "001000100000101000" => data <= "000000";
				when "001000100000101001" => data <= "000000";
				when "001000100000101010" => data <= "000000";
				when "001000100000101011" => data <= "000000";
				when "001000100000101100" => data <= "000000";
				when "001000100000101101" => data <= "000000";
				when "001000100000101110" => data <= "000000";
				when "001000100000101111" => data <= "000000";
				when "001000100000110000" => data <= "000000";
				when "001000100000110001" => data <= "000000";
				when "001000100000110010" => data <= "000000";
				when "001000100000110011" => data <= "000000";
				when "001000100000110100" => data <= "000000";
				when "001000100000110101" => data <= "000000";
				when "001000100000110110" => data <= "000000";
				when "001000100000110111" => data <= "000000";
				when "001000100000111000" => data <= "000000";
				when "001000100000111001" => data <= "000000";
				when "001000100000111010" => data <= "000000";
				when "001000100000111011" => data <= "000000";
				when "001000100000111100" => data <= "000000";
				when "001000100000111101" => data <= "000000";
				when "001000100000111110" => data <= "000000";
				when "001000100000111111" => data <= "000000";
				when "001000100001000000" => data <= "000000";
				when "001000100001000001" => data <= "000000";
				when "001000100001000010" => data <= "000000";
				when "001000100001000011" => data <= "000000";
				when "001000100001000100" => data <= "000000";
				when "001000100001000101" => data <= "000000";
				when "001000100001000110" => data <= "000000";
				when "001000100001000111" => data <= "000000";
				when "001000100001001000" => data <= "000000";
				when "001000100001001001" => data <= "000000";
				when "001000100001001010" => data <= "000000";
				when "001000100001001011" => data <= "000000";
				when "001000100001001100" => data <= "000000";
				when "001000100001001101" => data <= "000000";
				when "001000100001001110" => data <= "000000";
				when "001000100001001111" => data <= "000000";
				when "001000100001010000" => data <= "000000";
				when "001000100001010001" => data <= "000000";
				when "001000100001010010" => data <= "000000";
				when "001000100001010011" => data <= "000000";
				when "001000100001010100" => data <= "000000";
				when "001000100001010101" => data <= "000000";
				when "001000100001010110" => data <= "000000";
				when "001000100001010111" => data <= "000000";
				when "001000100001011000" => data <= "000000";
				when "001000100001011001" => data <= "000000";
				when "001000100001011010" => data <= "000000";
				when "001000100001011011" => data <= "000000";
				when "001000100001011100" => data <= "000000";
				when "001000100001011101" => data <= "000000";
				when "001000100001011110" => data <= "000000";
				when "001000100001011111" => data <= "000000";
				when "001000100001100000" => data <= "000000";
				when "001000100001100001" => data <= "000000";
				when "001000100001100010" => data <= "000000";
				when "001000100001100011" => data <= "000000";
				when "001000100001100100" => data <= "000000";
				when "001000100001100101" => data <= "000000";
				when "001000100001100110" => data <= "000000";
				when "001000100001100111" => data <= "000000";
				when "001000100001101000" => data <= "000000";
				when "001000100001101001" => data <= "000000";
				when "001000100001101010" => data <= "000000";
				when "001000100001101011" => data <= "000000";
				when "001000100001101100" => data <= "000000";
				when "001000100001101101" => data <= "000000";
				when "001000100001101110" => data <= "000000";
				when "001000100001101111" => data <= "000000";
				when "001000100001110000" => data <= "000000";
				when "001000100001110001" => data <= "000000";
				when "001000100001110010" => data <= "000000";
				when "001000100001110011" => data <= "000000";
				when "001000100001110100" => data <= "000000";
				when "001000100001110101" => data <= "000000";
				when "001000100001110110" => data <= "000000";
				when "001000100001110111" => data <= "000000";
				when "001000100001111000" => data <= "000000";
				when "001000100001111001" => data <= "000000";
				when "001000100001111010" => data <= "000000";
				when "001000100001111011" => data <= "000000";
				when "001000100001111100" => data <= "000000";
				when "001000100001111101" => data <= "000000";
				when "001000100001111110" => data <= "000000";
				when "001000100001111111" => data <= "000000";
				when "001000100010000000" => data <= "000000";
				when "001000100010000001" => data <= "000000";
				when "001000100010000010" => data <= "000000";
				when "001000100010000011" => data <= "000000";
				when "001000100010000100" => data <= "000000";
				when "001000100010000101" => data <= "000000";
				when "001000100010000110" => data <= "000000";
				when "001000100010000111" => data <= "000000";
				when "001000100010001000" => data <= "000000";
				when "001000100010001001" => data <= "000000";
				when "001000100010001010" => data <= "000000";
				when "001000100010001011" => data <= "000000";
				when "001000100010001100" => data <= "000000";
				when "001000100010001101" => data <= "000000";
				when "001000100010001110" => data <= "000000";
				when "001000100010001111" => data <= "000000";
				when "001000100010010000" => data <= "000000";
				when "001000100010010001" => data <= "000000";
				when "001000100010010010" => data <= "000000";
				when "001000100010010011" => data <= "000000";
				when "001000100010010100" => data <= "000000";
				when "001000100010010101" => data <= "000000";
				when "001000100010010110" => data <= "000000";
				when "001000100010010111" => data <= "000000";
				when "001000100010011000" => data <= "000000";
				when "001000100010011001" => data <= "000000";
				when "001000100010011010" => data <= "000000";
				when "001000100010011011" => data <= "000000";
				when "001000100010011100" => data <= "000000";
				when "001000100010011101" => data <= "000000";
				when "001000100010011110" => data <= "000000";
				when "001000100010011111" => data <= "000000";
				when "001000101000000000" => data <= "000000";
				when "001000101000000001" => data <= "000000";
				when "001000101000000010" => data <= "000000";
				when "001000101000000011" => data <= "000000";
				when "001000101000000100" => data <= "000000";
				when "001000101000000101" => data <= "000000";
				when "001000101000000110" => data <= "000000";
				when "001000101000000111" => data <= "000000";
				when "001000101000001000" => data <= "000000";
				when "001000101000001001" => data <= "000000";
				when "001000101000001010" => data <= "000000";
				when "001000101000001011" => data <= "000000";
				when "001000101000001100" => data <= "000000";
				when "001000101000001101" => data <= "000000";
				when "001000101000001110" => data <= "000000";
				when "001000101000001111" => data <= "000000";
				when "001000101000010000" => data <= "000000";
				when "001000101000010001" => data <= "000000";
				when "001000101000010010" => data <= "000000";
				when "001000101000010011" => data <= "000000";
				when "001000101000010100" => data <= "000000";
				when "001000101000010101" => data <= "000000";
				when "001000101000010110" => data <= "000000";
				when "001000101000010111" => data <= "000000";
				when "001000101000011000" => data <= "000000";
				when "001000101000011001" => data <= "000000";
				when "001000101000011010" => data <= "000000";
				when "001000101000011011" => data <= "000000";
				when "001000101000011100" => data <= "000000";
				when "001000101000011101" => data <= "000000";
				when "001000101000011110" => data <= "000000";
				when "001000101000011111" => data <= "000000";
				when "001000101000100000" => data <= "000000";
				when "001000101000100001" => data <= "000000";
				when "001000101000100010" => data <= "000000";
				when "001000101000100011" => data <= "000000";
				when "001000101000100100" => data <= "000000";
				when "001000101000100101" => data <= "000000";
				when "001000101000100110" => data <= "000000";
				when "001000101000100111" => data <= "000000";
				when "001000101000101000" => data <= "000000";
				when "001000101000101001" => data <= "000000";
				when "001000101000101010" => data <= "000000";
				when "001000101000101011" => data <= "000000";
				when "001000101000101100" => data <= "000000";
				when "001000101000101101" => data <= "000000";
				when "001000101000101110" => data <= "000000";
				when "001000101000101111" => data <= "000000";
				when "001000101000110000" => data <= "000000";
				when "001000101000110001" => data <= "000000";
				when "001000101000110010" => data <= "000000";
				when "001000101000110011" => data <= "000000";
				when "001000101000110100" => data <= "000000";
				when "001000101000110101" => data <= "000000";
				when "001000101000110110" => data <= "000000";
				when "001000101000110111" => data <= "000000";
				when "001000101000111000" => data <= "000000";
				when "001000101000111001" => data <= "000000";
				when "001000101000111010" => data <= "000000";
				when "001000101000111011" => data <= "000000";
				when "001000101000111100" => data <= "000000";
				when "001000101000111101" => data <= "000000";
				when "001000101000111110" => data <= "000000";
				when "001000101000111111" => data <= "000000";
				when "001000101001000000" => data <= "000000";
				when "001000101001000001" => data <= "000000";
				when "001000101001000010" => data <= "000000";
				when "001000101001000011" => data <= "000000";
				when "001000101001000100" => data <= "000000";
				when "001000101001000101" => data <= "000000";
				when "001000101001000110" => data <= "000000";
				when "001000101001000111" => data <= "000000";
				when "001000101001001000" => data <= "000000";
				when "001000101001001001" => data <= "000000";
				when "001000101001001010" => data <= "000000";
				when "001000101001001011" => data <= "000000";
				when "001000101001001100" => data <= "000000";
				when "001000101001001101" => data <= "000000";
				when "001000101001001110" => data <= "000000";
				when "001000101001001111" => data <= "000000";
				when "001000101001010000" => data <= "000000";
				when "001000101001010001" => data <= "000000";
				when "001000101001010010" => data <= "000000";
				when "001000101001010011" => data <= "000000";
				when "001000101001010100" => data <= "000000";
				when "001000101001010101" => data <= "000000";
				when "001000101001010110" => data <= "000000";
				when "001000101001010111" => data <= "000000";
				when "001000101001011000" => data <= "000000";
				when "001000101001011001" => data <= "000000";
				when "001000101001011010" => data <= "000000";
				when "001000101001011011" => data <= "000000";
				when "001000101001011100" => data <= "000000";
				when "001000101001011101" => data <= "000000";
				when "001000101001011110" => data <= "000000";
				when "001000101001011111" => data <= "000000";
				when "001000101001100000" => data <= "000000";
				when "001000101001100001" => data <= "000000";
				when "001000101001100010" => data <= "000000";
				when "001000101001100011" => data <= "000000";
				when "001000101001100100" => data <= "000000";
				when "001000101001100101" => data <= "000000";
				when "001000101001100110" => data <= "000000";
				when "001000101001100111" => data <= "000000";
				when "001000101001101000" => data <= "000000";
				when "001000101001101001" => data <= "000000";
				when "001000101001101010" => data <= "000000";
				when "001000101001101011" => data <= "000000";
				when "001000101001101100" => data <= "000000";
				when "001000101001101101" => data <= "000000";
				when "001000101001101110" => data <= "000000";
				when "001000101001101111" => data <= "000000";
				when "001000101001110000" => data <= "000000";
				when "001000101001110001" => data <= "000000";
				when "001000101001110010" => data <= "000000";
				when "001000101001110011" => data <= "000000";
				when "001000101001110100" => data <= "000000";
				when "001000101001110101" => data <= "000000";
				when "001000101001110110" => data <= "000000";
				when "001000101001110111" => data <= "000000";
				when "001000101001111000" => data <= "000000";
				when "001000101001111001" => data <= "000000";
				when "001000101001111010" => data <= "000000";
				when "001000101001111011" => data <= "000000";
				when "001000101001111100" => data <= "000000";
				when "001000101001111101" => data <= "000000";
				when "001000101001111110" => data <= "000000";
				when "001000101001111111" => data <= "000000";
				when "001000101010000000" => data <= "000000";
				when "001000101010000001" => data <= "000000";
				when "001000101010000010" => data <= "000000";
				when "001000101010000011" => data <= "000000";
				when "001000101010000100" => data <= "000000";
				when "001000101010000101" => data <= "000000";
				when "001000101010000110" => data <= "000000";
				when "001000101010000111" => data <= "000000";
				when "001000101010001000" => data <= "000000";
				when "001000101010001001" => data <= "000000";
				when "001000101010001010" => data <= "000000";
				when "001000101010001011" => data <= "000000";
				when "001000101010001100" => data <= "000000";
				when "001000101010001101" => data <= "000000";
				when "001000101010001110" => data <= "000000";
				when "001000101010001111" => data <= "000000";
				when "001000101010010000" => data <= "000000";
				when "001000101010010001" => data <= "000000";
				when "001000101010010010" => data <= "000000";
				when "001000101010010011" => data <= "000000";
				when "001000101010010100" => data <= "000000";
				when "001000101010010101" => data <= "000000";
				when "001000101010010110" => data <= "000000";
				when "001000101010010111" => data <= "000000";
				when "001000101010011000" => data <= "000000";
				when "001000101010011001" => data <= "000000";
				when "001000101010011010" => data <= "000000";
				when "001000101010011011" => data <= "000000";
				when "001000101010011100" => data <= "000000";
				when "001000101010011101" => data <= "000000";
				when "001000101010011110" => data <= "000000";
				when "001000101010011111" => data <= "000000";
				when "001000110000000000" => data <= "000000";
				when "001000110000000001" => data <= "000000";
				when "001000110000000010" => data <= "000000";
				when "001000110000000011" => data <= "000000";
				when "001000110000000100" => data <= "000000";
				when "001000110000000101" => data <= "000000";
				when "001000110000000110" => data <= "000000";
				when "001000110000000111" => data <= "000000";
				when "001000110000001000" => data <= "000000";
				when "001000110000001001" => data <= "000000";
				when "001000110000001010" => data <= "000000";
				when "001000110000001011" => data <= "000000";
				when "001000110000001100" => data <= "000000";
				when "001000110000001101" => data <= "000000";
				when "001000110000001110" => data <= "000000";
				when "001000110000001111" => data <= "000000";
				when "001000110000010000" => data <= "000000";
				when "001000110000010001" => data <= "000000";
				when "001000110000010010" => data <= "000000";
				when "001000110000010011" => data <= "000000";
				when "001000110000010100" => data <= "000000";
				when "001000110000010101" => data <= "000000";
				when "001000110000010110" => data <= "000000";
				when "001000110000010111" => data <= "000000";
				when "001000110000011000" => data <= "000000";
				when "001000110000011001" => data <= "000000";
				when "001000110000011010" => data <= "000000";
				when "001000110000011011" => data <= "000000";
				when "001000110000011100" => data <= "000000";
				when "001000110000011101" => data <= "000000";
				when "001000110000011110" => data <= "000000";
				when "001000110000011111" => data <= "000000";
				when "001000110000100000" => data <= "000000";
				when "001000110000100001" => data <= "000000";
				when "001000110000100010" => data <= "000000";
				when "001000110000100011" => data <= "000000";
				when "001000110000100100" => data <= "000000";
				when "001000110000100101" => data <= "000000";
				when "001000110000100110" => data <= "000000";
				when "001000110000100111" => data <= "000000";
				when "001000110000101000" => data <= "000000";
				when "001000110000101001" => data <= "000000";
				when "001000110000101010" => data <= "000000";
				when "001000110000101011" => data <= "000000";
				when "001000110000101100" => data <= "000000";
				when "001000110000101101" => data <= "000000";
				when "001000110000101110" => data <= "000000";
				when "001000110000101111" => data <= "000000";
				when "001000110000110000" => data <= "000000";
				when "001000110000110001" => data <= "000000";
				when "001000110000110010" => data <= "000000";
				when "001000110000110011" => data <= "000000";
				when "001000110000110100" => data <= "000000";
				when "001000110000110101" => data <= "000000";
				when "001000110000110110" => data <= "000000";
				when "001000110000110111" => data <= "000000";
				when "001000110000111000" => data <= "000000";
				when "001000110000111001" => data <= "000000";
				when "001000110000111010" => data <= "000000";
				when "001000110000111011" => data <= "000000";
				when "001000110000111100" => data <= "000000";
				when "001000110000111101" => data <= "000000";
				when "001000110000111110" => data <= "000000";
				when "001000110000111111" => data <= "000000";
				when "001000110001000000" => data <= "000000";
				when "001000110001000001" => data <= "000000";
				when "001000110001000010" => data <= "000000";
				when "001000110001000011" => data <= "000000";
				when "001000110001000100" => data <= "000000";
				when "001000110001000101" => data <= "000000";
				when "001000110001000110" => data <= "000000";
				when "001000110001000111" => data <= "000000";
				when "001000110001001000" => data <= "000000";
				when "001000110001001001" => data <= "000000";
				when "001000110001001010" => data <= "000000";
				when "001000110001001011" => data <= "000000";
				when "001000110001001100" => data <= "000000";
				when "001000110001001101" => data <= "000000";
				when "001000110001001110" => data <= "000000";
				when "001000110001001111" => data <= "000000";
				when "001000110001010000" => data <= "000000";
				when "001000110001010001" => data <= "000000";
				when "001000110001010010" => data <= "000000";
				when "001000110001010011" => data <= "000000";
				when "001000110001010100" => data <= "000000";
				when "001000110001010101" => data <= "000000";
				when "001000110001010110" => data <= "000000";
				when "001000110001010111" => data <= "000000";
				when "001000110001011000" => data <= "000000";
				when "001000110001011001" => data <= "000000";
				when "001000110001011010" => data <= "000000";
				when "001000110001011011" => data <= "000000";
				when "001000110001011100" => data <= "000000";
				when "001000110001011101" => data <= "000000";
				when "001000110001011110" => data <= "000000";
				when "001000110001011111" => data <= "000000";
				when "001000110001100000" => data <= "000000";
				when "001000110001100001" => data <= "000000";
				when "001000110001100010" => data <= "000000";
				when "001000110001100011" => data <= "000000";
				when "001000110001100100" => data <= "000000";
				when "001000110001100101" => data <= "000000";
				when "001000110001100110" => data <= "000000";
				when "001000110001100111" => data <= "000000";
				when "001000110001101000" => data <= "000000";
				when "001000110001101001" => data <= "000000";
				when "001000110001101010" => data <= "000000";
				when "001000110001101011" => data <= "000000";
				when "001000110001101100" => data <= "000000";
				when "001000110001101101" => data <= "000000";
				when "001000110001101110" => data <= "000000";
				when "001000110001101111" => data <= "000000";
				when "001000110001110000" => data <= "000000";
				when "001000110001110001" => data <= "000000";
				when "001000110001110010" => data <= "000000";
				when "001000110001110011" => data <= "000000";
				when "001000110001110100" => data <= "000000";
				when "001000110001110101" => data <= "000000";
				when "001000110001110110" => data <= "000000";
				when "001000110001110111" => data <= "000000";
				when "001000110001111000" => data <= "000000";
				when "001000110001111001" => data <= "000000";
				when "001000110001111010" => data <= "000000";
				when "001000110001111011" => data <= "000000";
				when "001000110001111100" => data <= "000000";
				when "001000110001111101" => data <= "000000";
				when "001000110001111110" => data <= "000000";
				when "001000110001111111" => data <= "000000";
				when "001000110010000000" => data <= "000000";
				when "001000110010000001" => data <= "000000";
				when "001000110010000010" => data <= "000000";
				when "001000110010000011" => data <= "000000";
				when "001000110010000100" => data <= "000000";
				when "001000110010000101" => data <= "000000";
				when "001000110010000110" => data <= "000000";
				when "001000110010000111" => data <= "000000";
				when "001000110010001000" => data <= "000000";
				when "001000110010001001" => data <= "000000";
				when "001000110010001010" => data <= "000000";
				when "001000110010001011" => data <= "000000";
				when "001000110010001100" => data <= "000000";
				when "001000110010001101" => data <= "000000";
				when "001000110010001110" => data <= "000000";
				when "001000110010001111" => data <= "000000";
				when "001000110010010000" => data <= "000000";
				when "001000110010010001" => data <= "000000";
				when "001000110010010010" => data <= "000000";
				when "001000110010010011" => data <= "000000";
				when "001000110010010100" => data <= "000000";
				when "001000110010010101" => data <= "000000";
				when "001000110010010110" => data <= "000000";
				when "001000110010010111" => data <= "000000";
				when "001000110010011000" => data <= "000000";
				when "001000110010011001" => data <= "000000";
				when "001000110010011010" => data <= "000000";
				when "001000110010011011" => data <= "000000";
				when "001000110010011100" => data <= "000000";
				when "001000110010011101" => data <= "000000";
				when "001000110010011110" => data <= "000000";
				when "001000110010011111" => data <= "000000";
				when "001000111000000000" => data <= "000000";
				when "001000111000000001" => data <= "000000";
				when "001000111000000010" => data <= "000000";
				when "001000111000000011" => data <= "000000";
				when "001000111000000100" => data <= "000000";
				when "001000111000000101" => data <= "000000";
				when "001000111000000110" => data <= "000000";
				when "001000111000000111" => data <= "000000";
				when "001000111000001000" => data <= "000000";
				when "001000111000001001" => data <= "000000";
				when "001000111000001010" => data <= "000000";
				when "001000111000001011" => data <= "000000";
				when "001000111000001100" => data <= "000000";
				when "001000111000001101" => data <= "000000";
				when "001000111000001110" => data <= "000000";
				when "001000111000001111" => data <= "000000";
				when "001000111000010000" => data <= "000000";
				when "001000111000010001" => data <= "000000";
				when "001000111000010010" => data <= "000000";
				when "001000111000010011" => data <= "000000";
				when "001000111000010100" => data <= "000000";
				when "001000111000010101" => data <= "000000";
				when "001000111000010110" => data <= "000000";
				when "001000111000010111" => data <= "000000";
				when "001000111000011000" => data <= "000000";
				when "001000111000011001" => data <= "000000";
				when "001000111000011010" => data <= "000000";
				when "001000111000011011" => data <= "000000";
				when "001000111000011100" => data <= "000000";
				when "001000111000011101" => data <= "000000";
				when "001000111000011110" => data <= "000000";
				when "001000111000011111" => data <= "000000";
				when "001000111000100000" => data <= "000000";
				when "001000111000100001" => data <= "000000";
				when "001000111000100010" => data <= "000000";
				when "001000111000100011" => data <= "000000";
				when "001000111000100100" => data <= "000000";
				when "001000111000100101" => data <= "000000";
				when "001000111000100110" => data <= "000000";
				when "001000111000100111" => data <= "000000";
				when "001000111000101000" => data <= "000000";
				when "001000111000101001" => data <= "000000";
				when "001000111000101010" => data <= "000000";
				when "001000111000101011" => data <= "000000";
				when "001000111000101100" => data <= "000000";
				when "001000111000101101" => data <= "000000";
				when "001000111000101110" => data <= "000000";
				when "001000111000101111" => data <= "000000";
				when "001000111000110000" => data <= "000000";
				when "001000111000110001" => data <= "000000";
				when "001000111000110010" => data <= "000000";
				when "001000111000110011" => data <= "000000";
				when "001000111000110100" => data <= "000000";
				when "001000111000110101" => data <= "000000";
				when "001000111000110110" => data <= "000000";
				when "001000111000110111" => data <= "000000";
				when "001000111000111000" => data <= "000000";
				when "001000111000111001" => data <= "000000";
				when "001000111000111010" => data <= "000000";
				when "001000111000111011" => data <= "000000";
				when "001000111000111100" => data <= "000000";
				when "001000111000111101" => data <= "000000";
				when "001000111000111110" => data <= "000000";
				when "001000111000111111" => data <= "000000";
				when "001000111001000000" => data <= "000000";
				when "001000111001000001" => data <= "000000";
				when "001000111001000010" => data <= "000000";
				when "001000111001000011" => data <= "000000";
				when "001000111001000100" => data <= "000000";
				when "001000111001000101" => data <= "000000";
				when "001000111001000110" => data <= "000000";
				when "001000111001000111" => data <= "000000";
				when "001000111001001000" => data <= "000000";
				when "001000111001001001" => data <= "000000";
				when "001000111001001010" => data <= "000000";
				when "001000111001001011" => data <= "000000";
				when "001000111001001100" => data <= "000000";
				when "001000111001001101" => data <= "000000";
				when "001000111001001110" => data <= "000000";
				when "001000111001001111" => data <= "000000";
				when "001000111001010000" => data <= "000000";
				when "001000111001010001" => data <= "000000";
				when "001000111001010010" => data <= "000000";
				when "001000111001010011" => data <= "000000";
				when "001000111001010100" => data <= "000000";
				when "001000111001010101" => data <= "000000";
				when "001000111001010110" => data <= "000000";
				when "001000111001010111" => data <= "000000";
				when "001000111001011000" => data <= "000000";
				when "001000111001011001" => data <= "000000";
				when "001000111001011010" => data <= "000000";
				when "001000111001011011" => data <= "000000";
				when "001000111001011100" => data <= "000000";
				when "001000111001011101" => data <= "000000";
				when "001000111001011110" => data <= "000000";
				when "001000111001011111" => data <= "000000";
				when "001000111001100000" => data <= "000000";
				when "001000111001100001" => data <= "000000";
				when "001000111001100010" => data <= "000000";
				when "001000111001100011" => data <= "000000";
				when "001000111001100100" => data <= "000000";
				when "001000111001100101" => data <= "000000";
				when "001000111001100110" => data <= "000000";
				when "001000111001100111" => data <= "000000";
				when "001000111001101000" => data <= "000000";
				when "001000111001101001" => data <= "000000";
				when "001000111001101010" => data <= "000000";
				when "001000111001101011" => data <= "000000";
				when "001000111001101100" => data <= "000000";
				when "001000111001101101" => data <= "000000";
				when "001000111001101110" => data <= "000000";
				when "001000111001101111" => data <= "000000";
				when "001000111001110000" => data <= "000000";
				when "001000111001110001" => data <= "000000";
				when "001000111001110010" => data <= "000000";
				when "001000111001110011" => data <= "000000";
				when "001000111001110100" => data <= "000000";
				when "001000111001110101" => data <= "000000";
				when "001000111001110110" => data <= "000000";
				when "001000111001110111" => data <= "000000";
				when "001000111001111000" => data <= "000000";
				when "001000111001111001" => data <= "000000";
				when "001000111001111010" => data <= "000000";
				when "001000111001111011" => data <= "000000";
				when "001000111001111100" => data <= "000000";
				when "001000111001111101" => data <= "000000";
				when "001000111001111110" => data <= "000000";
				when "001000111001111111" => data <= "000000";
				when "001000111010000000" => data <= "000000";
				when "001000111010000001" => data <= "000000";
				when "001000111010000010" => data <= "000000";
				when "001000111010000011" => data <= "000000";
				when "001000111010000100" => data <= "000000";
				when "001000111010000101" => data <= "000000";
				when "001000111010000110" => data <= "000000";
				when "001000111010000111" => data <= "000000";
				when "001000111010001000" => data <= "000000";
				when "001000111010001001" => data <= "000000";
				when "001000111010001010" => data <= "000000";
				when "001000111010001011" => data <= "000000";
				when "001000111010001100" => data <= "000000";
				when "001000111010001101" => data <= "000000";
				when "001000111010001110" => data <= "000000";
				when "001000111010001111" => data <= "000000";
				when "001000111010010000" => data <= "000000";
				when "001000111010010001" => data <= "000000";
				when "001000111010010010" => data <= "000000";
				when "001000111010010011" => data <= "000000";
				when "001000111010010100" => data <= "000000";
				when "001000111010010101" => data <= "000000";
				when "001000111010010110" => data <= "000000";
				when "001000111010010111" => data <= "000000";
				when "001000111010011000" => data <= "000000";
				when "001000111010011001" => data <= "000000";
				when "001000111010011010" => data <= "000000";
				when "001000111010011011" => data <= "000000";
				when "001000111010011100" => data <= "000000";
				when "001000111010011101" => data <= "000000";
				when "001000111010011110" => data <= "000000";
				when "001000111010011111" => data <= "000000";
				when "001001000000000000" => data <= "000000";
				when "001001000000000001" => data <= "000000";
				when "001001000000000010" => data <= "000000";
				when "001001000000000011" => data <= "000000";
				when "001001000000000100" => data <= "000000";
				when "001001000000000101" => data <= "000000";
				when "001001000000000110" => data <= "000000";
				when "001001000000000111" => data <= "000000";
				when "001001000000001000" => data <= "000000";
				when "001001000000001001" => data <= "000000";
				when "001001000000001010" => data <= "000000";
				when "001001000000001011" => data <= "000000";
				when "001001000000001100" => data <= "000000";
				when "001001000000001101" => data <= "000000";
				when "001001000000001110" => data <= "000000";
				when "001001000000001111" => data <= "000000";
				when "001001000000010000" => data <= "000000";
				when "001001000000010001" => data <= "000000";
				when "001001000000010010" => data <= "000000";
				when "001001000000010011" => data <= "000000";
				when "001001000000010100" => data <= "000000";
				when "001001000000010101" => data <= "000000";
				when "001001000000010110" => data <= "000000";
				when "001001000000010111" => data <= "000000";
				when "001001000000011000" => data <= "000000";
				when "001001000000011001" => data <= "000000";
				when "001001000000011010" => data <= "000000";
				when "001001000000011011" => data <= "000000";
				when "001001000000011100" => data <= "000000";
				when "001001000000011101" => data <= "000000";
				when "001001000000011110" => data <= "000000";
				when "001001000000011111" => data <= "000000";
				when "001001000000100000" => data <= "000000";
				when "001001000000100001" => data <= "000000";
				when "001001000000100010" => data <= "000000";
				when "001001000000100011" => data <= "000000";
				when "001001000000100100" => data <= "000000";
				when "001001000000100101" => data <= "000000";
				when "001001000000100110" => data <= "000000";
				when "001001000000100111" => data <= "000000";
				when "001001000000101000" => data <= "000000";
				when "001001000000101001" => data <= "000000";
				when "001001000000101010" => data <= "000000";
				when "001001000000101011" => data <= "000000";
				when "001001000000101100" => data <= "000000";
				when "001001000000101101" => data <= "000000";
				when "001001000000101110" => data <= "000000";
				when "001001000000101111" => data <= "000000";
				when "001001000000110000" => data <= "000000";
				when "001001000000110001" => data <= "000000";
				when "001001000000110010" => data <= "000000";
				when "001001000000110011" => data <= "000000";
				when "001001000000110100" => data <= "000000";
				when "001001000000110101" => data <= "000000";
				when "001001000000110110" => data <= "000000";
				when "001001000000110111" => data <= "000000";
				when "001001000000111000" => data <= "000000";
				when "001001000000111001" => data <= "000000";
				when "001001000000111010" => data <= "000000";
				when "001001000000111011" => data <= "000000";
				when "001001000000111100" => data <= "000000";
				when "001001000000111101" => data <= "000000";
				when "001001000000111110" => data <= "000000";
				when "001001000000111111" => data <= "000000";
				when "001001000001000000" => data <= "000000";
				when "001001000001000001" => data <= "000000";
				when "001001000001000010" => data <= "000000";
				when "001001000001000011" => data <= "000000";
				when "001001000001000100" => data <= "000000";
				when "001001000001000101" => data <= "000000";
				when "001001000001000110" => data <= "000000";
				when "001001000001000111" => data <= "000000";
				when "001001000001001000" => data <= "000000";
				when "001001000001001001" => data <= "000000";
				when "001001000001001010" => data <= "000000";
				when "001001000001001011" => data <= "000000";
				when "001001000001001100" => data <= "000000";
				when "001001000001001101" => data <= "000000";
				when "001001000001001110" => data <= "000000";
				when "001001000001001111" => data <= "000000";
				when "001001000001010000" => data <= "000000";
				when "001001000001010001" => data <= "000000";
				when "001001000001010010" => data <= "000000";
				when "001001000001010011" => data <= "000000";
				when "001001000001010100" => data <= "000000";
				when "001001000001010101" => data <= "000000";
				when "001001000001010110" => data <= "000000";
				when "001001000001010111" => data <= "000000";
				when "001001000001011000" => data <= "000000";
				when "001001000001011001" => data <= "000000";
				when "001001000001011010" => data <= "000000";
				when "001001000001011011" => data <= "000000";
				when "001001000001011100" => data <= "000000";
				when "001001000001011101" => data <= "000000";
				when "001001000001011110" => data <= "000000";
				when "001001000001011111" => data <= "000000";
				when "001001000001100000" => data <= "000000";
				when "001001000001100001" => data <= "000000";
				when "001001000001100010" => data <= "000000";
				when "001001000001100011" => data <= "000000";
				when "001001000001100100" => data <= "000000";
				when "001001000001100101" => data <= "000000";
				when "001001000001100110" => data <= "000000";
				when "001001000001100111" => data <= "000000";
				when "001001000001101000" => data <= "000000";
				when "001001000001101001" => data <= "000000";
				when "001001000001101010" => data <= "000000";
				when "001001000001101011" => data <= "000000";
				when "001001000001101100" => data <= "000000";
				when "001001000001101101" => data <= "000000";
				when "001001000001101110" => data <= "000000";
				when "001001000001101111" => data <= "000000";
				when "001001000001110000" => data <= "000000";
				when "001001000001110001" => data <= "000000";
				when "001001000001110010" => data <= "000000";
				when "001001000001110011" => data <= "000000";
				when "001001000001110100" => data <= "000000";
				when "001001000001110101" => data <= "000000";
				when "001001000001110110" => data <= "000000";
				when "001001000001110111" => data <= "000000";
				when "001001000001111000" => data <= "000000";
				when "001001000001111001" => data <= "000000";
				when "001001000001111010" => data <= "000000";
				when "001001000001111011" => data <= "000000";
				when "001001000001111100" => data <= "000000";
				when "001001000001111101" => data <= "000000";
				when "001001000001111110" => data <= "000000";
				when "001001000001111111" => data <= "000000";
				when "001001000010000000" => data <= "000000";
				when "001001000010000001" => data <= "000000";
				when "001001000010000010" => data <= "000000";
				when "001001000010000011" => data <= "000000";
				when "001001000010000100" => data <= "000000";
				when "001001000010000101" => data <= "000000";
				when "001001000010000110" => data <= "000000";
				when "001001000010000111" => data <= "000000";
				when "001001000010001000" => data <= "000000";
				when "001001000010001001" => data <= "000000";
				when "001001000010001010" => data <= "000000";
				when "001001000010001011" => data <= "000000";
				when "001001000010001100" => data <= "000000";
				when "001001000010001101" => data <= "000000";
				when "001001000010001110" => data <= "000000";
				when "001001000010001111" => data <= "000000";
				when "001001000010010000" => data <= "000000";
				when "001001000010010001" => data <= "000000";
				when "001001000010010010" => data <= "000000";
				when "001001000010010011" => data <= "000000";
				when "001001000010010100" => data <= "000000";
				when "001001000010010101" => data <= "000000";
				when "001001000010010110" => data <= "000000";
				when "001001000010010111" => data <= "000000";
				when "001001000010011000" => data <= "000000";
				when "001001000010011001" => data <= "000000";
				when "001001000010011010" => data <= "000000";
				when "001001000010011011" => data <= "000000";
				when "001001000010011100" => data <= "000000";
				when "001001000010011101" => data <= "000000";
				when "001001000010011110" => data <= "000000";
				when "001001000010011111" => data <= "000000";
				when "001001001000000000" => data <= "000000";
				when "001001001000000001" => data <= "000000";
				when "001001001000000010" => data <= "000000";
				when "001001001000000011" => data <= "000000";
				when "001001001000000100" => data <= "000000";
				when "001001001000000101" => data <= "000000";
				when "001001001000000110" => data <= "000000";
				when "001001001000000111" => data <= "000000";
				when "001001001000001000" => data <= "000000";
				when "001001001000001001" => data <= "000000";
				when "001001001000001010" => data <= "000000";
				when "001001001000001011" => data <= "000000";
				when "001001001000001100" => data <= "000000";
				when "001001001000001101" => data <= "000000";
				when "001001001000001110" => data <= "000000";
				when "001001001000001111" => data <= "000000";
				when "001001001000010000" => data <= "000000";
				when "001001001000010001" => data <= "000000";
				when "001001001000010010" => data <= "000000";
				when "001001001000010011" => data <= "000000";
				when "001001001000010100" => data <= "000000";
				when "001001001000010101" => data <= "000000";
				when "001001001000010110" => data <= "000000";
				when "001001001000010111" => data <= "000000";
				when "001001001000011000" => data <= "000000";
				when "001001001000011001" => data <= "000000";
				when "001001001000011010" => data <= "000000";
				when "001001001000011011" => data <= "000000";
				when "001001001000011100" => data <= "000000";
				when "001001001000011101" => data <= "000000";
				when "001001001000011110" => data <= "000000";
				when "001001001000011111" => data <= "000000";
				when "001001001000100000" => data <= "000000";
				when "001001001000100001" => data <= "000000";
				when "001001001000100010" => data <= "000000";
				when "001001001000100011" => data <= "000000";
				when "001001001000100100" => data <= "000000";
				when "001001001000100101" => data <= "000000";
				when "001001001000100110" => data <= "000000";
				when "001001001000100111" => data <= "000000";
				when "001001001000101000" => data <= "000000";
				when "001001001000101001" => data <= "000000";
				when "001001001000101010" => data <= "000000";
				when "001001001000101011" => data <= "000000";
				when "001001001000101100" => data <= "000000";
				when "001001001000101101" => data <= "000000";
				when "001001001000101110" => data <= "000000";
				when "001001001000101111" => data <= "000000";
				when "001001001000110000" => data <= "000000";
				when "001001001000110001" => data <= "000000";
				when "001001001000110010" => data <= "000000";
				when "001001001000110011" => data <= "000000";
				when "001001001000110100" => data <= "000000";
				when "001001001000110101" => data <= "000000";
				when "001001001000110110" => data <= "000000";
				when "001001001000110111" => data <= "000000";
				when "001001001000111000" => data <= "000000";
				when "001001001000111001" => data <= "000000";
				when "001001001000111010" => data <= "000000";
				when "001001001000111011" => data <= "000000";
				when "001001001000111100" => data <= "000000";
				when "001001001000111101" => data <= "000000";
				when "001001001000111110" => data <= "000000";
				when "001001001000111111" => data <= "000000";
				when "001001001001000000" => data <= "000000";
				when "001001001001000001" => data <= "000000";
				when "001001001001000010" => data <= "000000";
				when "001001001001000011" => data <= "000000";
				when "001001001001000100" => data <= "000000";
				when "001001001001000101" => data <= "000000";
				when "001001001001000110" => data <= "000000";
				when "001001001001000111" => data <= "000000";
				when "001001001001001000" => data <= "000000";
				when "001001001001001001" => data <= "000000";
				when "001001001001001010" => data <= "000000";
				when "001001001001001011" => data <= "000000";
				when "001001001001001100" => data <= "000000";
				when "001001001001001101" => data <= "000000";
				when "001001001001001110" => data <= "000000";
				when "001001001001001111" => data <= "000000";
				when "001001001001010000" => data <= "000000";
				when "001001001001010001" => data <= "000000";
				when "001001001001010010" => data <= "000000";
				when "001001001001010011" => data <= "000000";
				when "001001001001010100" => data <= "000000";
				when "001001001001010101" => data <= "000000";
				when "001001001001010110" => data <= "000000";
				when "001001001001010111" => data <= "000000";
				when "001001001001011000" => data <= "000000";
				when "001001001001011001" => data <= "000000";
				when "001001001001011010" => data <= "000000";
				when "001001001001011011" => data <= "000000";
				when "001001001001011100" => data <= "000000";
				when "001001001001011101" => data <= "000000";
				when "001001001001011110" => data <= "000000";
				when "001001001001011111" => data <= "000000";
				when "001001001001100000" => data <= "000000";
				when "001001001001100001" => data <= "000000";
				when "001001001001100010" => data <= "000000";
				when "001001001001100011" => data <= "000000";
				when "001001001001100100" => data <= "000000";
				when "001001001001100101" => data <= "000000";
				when "001001001001100110" => data <= "000000";
				when "001001001001100111" => data <= "000000";
				when "001001001001101000" => data <= "000000";
				when "001001001001101001" => data <= "000000";
				when "001001001001101010" => data <= "000000";
				when "001001001001101011" => data <= "000000";
				when "001001001001101100" => data <= "000000";
				when "001001001001101101" => data <= "000000";
				when "001001001001101110" => data <= "000000";
				when "001001001001101111" => data <= "000000";
				when "001001001001110000" => data <= "000000";
				when "001001001001110001" => data <= "000000";
				when "001001001001110010" => data <= "000000";
				when "001001001001110011" => data <= "000000";
				when "001001001001110100" => data <= "000000";
				when "001001001001110101" => data <= "000000";
				when "001001001001110110" => data <= "000000";
				when "001001001001110111" => data <= "000000";
				when "001001001001111000" => data <= "000000";
				when "001001001001111001" => data <= "000000";
				when "001001001001111010" => data <= "000000";
				when "001001001001111011" => data <= "000000";
				when "001001001001111100" => data <= "000000";
				when "001001001001111101" => data <= "000000";
				when "001001001001111110" => data <= "000000";
				when "001001001001111111" => data <= "000000";
				when "001001001010000000" => data <= "000000";
				when "001001001010000001" => data <= "000000";
				when "001001001010000010" => data <= "000000";
				when "001001001010000011" => data <= "000000";
				when "001001001010000100" => data <= "000000";
				when "001001001010000101" => data <= "000000";
				when "001001001010000110" => data <= "000000";
				when "001001001010000111" => data <= "000000";
				when "001001001010001000" => data <= "000000";
				when "001001001010001001" => data <= "000000";
				when "001001001010001010" => data <= "000000";
				when "001001001010001011" => data <= "000000";
				when "001001001010001100" => data <= "000000";
				when "001001001010001101" => data <= "000000";
				when "001001001010001110" => data <= "000000";
				when "001001001010001111" => data <= "000000";
				when "001001001010010000" => data <= "000000";
				when "001001001010010001" => data <= "000000";
				when "001001001010010010" => data <= "000000";
				when "001001001010010011" => data <= "000000";
				when "001001001010010100" => data <= "000000";
				when "001001001010010101" => data <= "000000";
				when "001001001010010110" => data <= "000000";
				when "001001001010010111" => data <= "000000";
				when "001001001010011000" => data <= "000000";
				when "001001001010011001" => data <= "000000";
				when "001001001010011010" => data <= "000000";
				when "001001001010011011" => data <= "000000";
				when "001001001010011100" => data <= "000000";
				when "001001001010011101" => data <= "000000";
				when "001001001010011110" => data <= "000000";
				when "001001001010011111" => data <= "000000";
				when "001001010000000000" => data <= "000000";
				when "001001010000000001" => data <= "000000";
				when "001001010000000010" => data <= "000000";
				when "001001010000000011" => data <= "000000";
				when "001001010000000100" => data <= "000000";
				when "001001010000000101" => data <= "000000";
				when "001001010000000110" => data <= "000000";
				when "001001010000000111" => data <= "000000";
				when "001001010000001000" => data <= "000000";
				when "001001010000001001" => data <= "000000";
				when "001001010000001010" => data <= "000000";
				when "001001010000001011" => data <= "000000";
				when "001001010000001100" => data <= "000000";
				when "001001010000001101" => data <= "000000";
				when "001001010000001110" => data <= "000000";
				when "001001010000001111" => data <= "000000";
				when "001001010000010000" => data <= "000000";
				when "001001010000010001" => data <= "000000";
				when "001001010000010010" => data <= "000000";
				when "001001010000010011" => data <= "000000";
				when "001001010000010100" => data <= "000000";
				when "001001010000010101" => data <= "000000";
				when "001001010000010110" => data <= "000000";
				when "001001010000010111" => data <= "000000";
				when "001001010000011000" => data <= "000000";
				when "001001010000011001" => data <= "000000";
				when "001001010000011010" => data <= "000000";
				when "001001010000011011" => data <= "000000";
				when "001001010000011100" => data <= "000000";
				when "001001010000011101" => data <= "000000";
				when "001001010000011110" => data <= "000000";
				when "001001010000011111" => data <= "000000";
				when "001001010000100000" => data <= "000000";
				when "001001010000100001" => data <= "000000";
				when "001001010000100010" => data <= "000000";
				when "001001010000100011" => data <= "000000";
				when "001001010000100100" => data <= "000000";
				when "001001010000100101" => data <= "000000";
				when "001001010000100110" => data <= "000000";
				when "001001010000100111" => data <= "000000";
				when "001001010000101000" => data <= "000000";
				when "001001010000101001" => data <= "000000";
				when "001001010000101010" => data <= "000000";
				when "001001010000101011" => data <= "000000";
				when "001001010000101100" => data <= "000000";
				when "001001010000101101" => data <= "000000";
				when "001001010000101110" => data <= "000000";
				when "001001010000101111" => data <= "000000";
				when "001001010000110000" => data <= "000000";
				when "001001010000110001" => data <= "000000";
				when "001001010000110010" => data <= "000000";
				when "001001010000110011" => data <= "000000";
				when "001001010000110100" => data <= "000000";
				when "001001010000110101" => data <= "000000";
				when "001001010000110110" => data <= "000000";
				when "001001010000110111" => data <= "000000";
				when "001001010000111000" => data <= "000000";
				when "001001010000111001" => data <= "000000";
				when "001001010000111010" => data <= "000000";
				when "001001010000111011" => data <= "000000";
				when "001001010000111100" => data <= "000000";
				when "001001010000111101" => data <= "000000";
				when "001001010000111110" => data <= "000000";
				when "001001010000111111" => data <= "000000";
				when "001001010001000000" => data <= "000000";
				when "001001010001000001" => data <= "000000";
				when "001001010001000010" => data <= "000000";
				when "001001010001000011" => data <= "000000";
				when "001001010001000100" => data <= "000000";
				when "001001010001000101" => data <= "000000";
				when "001001010001000110" => data <= "000000";
				when "001001010001000111" => data <= "000000";
				when "001001010001001000" => data <= "000000";
				when "001001010001001001" => data <= "000000";
				when "001001010001001010" => data <= "000000";
				when "001001010001001011" => data <= "000000";
				when "001001010001001100" => data <= "000000";
				when "001001010001001101" => data <= "000000";
				when "001001010001001110" => data <= "000000";
				when "001001010001001111" => data <= "000000";
				when "001001010001010000" => data <= "000000";
				when "001001010001010001" => data <= "000000";
				when "001001010001010010" => data <= "000000";
				when "001001010001010011" => data <= "000000";
				when "001001010001010100" => data <= "000000";
				when "001001010001010101" => data <= "000000";
				when "001001010001010110" => data <= "000000";
				when "001001010001010111" => data <= "000000";
				when "001001010001011000" => data <= "000000";
				when "001001010001011001" => data <= "000000";
				when "001001010001011010" => data <= "000000";
				when "001001010001011011" => data <= "000000";
				when "001001010001011100" => data <= "000000";
				when "001001010001011101" => data <= "000000";
				when "001001010001011110" => data <= "000000";
				when "001001010001011111" => data <= "000000";
				when "001001010001100000" => data <= "000000";
				when "001001010001100001" => data <= "000000";
				when "001001010001100010" => data <= "000000";
				when "001001010001100011" => data <= "000000";
				when "001001010001100100" => data <= "000000";
				when "001001010001100101" => data <= "000000";
				when "001001010001100110" => data <= "000000";
				when "001001010001100111" => data <= "000000";
				when "001001010001101000" => data <= "000000";
				when "001001010001101001" => data <= "000000";
				when "001001010001101010" => data <= "000000";
				when "001001010001101011" => data <= "000000";
				when "001001010001101100" => data <= "000000";
				when "001001010001101101" => data <= "000000";
				when "001001010001101110" => data <= "000000";
				when "001001010001101111" => data <= "000000";
				when "001001010001110000" => data <= "000000";
				when "001001010001110001" => data <= "000000";
				when "001001010001110010" => data <= "000000";
				when "001001010001110011" => data <= "000000";
				when "001001010001110100" => data <= "000000";
				when "001001010001110101" => data <= "000000";
				when "001001010001110110" => data <= "000000";
				when "001001010001110111" => data <= "000000";
				when "001001010001111000" => data <= "000000";
				when "001001010001111001" => data <= "000000";
				when "001001010001111010" => data <= "000000";
				when "001001010001111011" => data <= "000000";
				when "001001010001111100" => data <= "000000";
				when "001001010001111101" => data <= "000000";
				when "001001010001111110" => data <= "000000";
				when "001001010001111111" => data <= "000000";
				when "001001010010000000" => data <= "000000";
				when "001001010010000001" => data <= "000000";
				when "001001010010000010" => data <= "000000";
				when "001001010010000011" => data <= "000000";
				when "001001010010000100" => data <= "000000";
				when "001001010010000101" => data <= "000000";
				when "001001010010000110" => data <= "000000";
				when "001001010010000111" => data <= "000000";
				when "001001010010001000" => data <= "000000";
				when "001001010010001001" => data <= "000000";
				when "001001010010001010" => data <= "000000";
				when "001001010010001011" => data <= "000000";
				when "001001010010001100" => data <= "000000";
				when "001001010010001101" => data <= "000000";
				when "001001010010001110" => data <= "000000";
				when "001001010010001111" => data <= "000000";
				when "001001010010010000" => data <= "000000";
				when "001001010010010001" => data <= "000000";
				when "001001010010010010" => data <= "000000";
				when "001001010010010011" => data <= "000000";
				when "001001010010010100" => data <= "000000";
				when "001001010010010101" => data <= "000000";
				when "001001010010010110" => data <= "000000";
				when "001001010010010111" => data <= "000000";
				when "001001010010011000" => data <= "000000";
				when "001001010010011001" => data <= "000000";
				when "001001010010011010" => data <= "000000";
				when "001001010010011011" => data <= "000000";
				when "001001010010011100" => data <= "000000";
				when "001001010010011101" => data <= "000000";
				when "001001010010011110" => data <= "000000";
				when "001001010010011111" => data <= "000000";
				when "001001011000000000" => data <= "000000";
				when "001001011000000001" => data <= "000000";
				when "001001011000000010" => data <= "000000";
				when "001001011000000011" => data <= "000000";
				when "001001011000000100" => data <= "000000";
				when "001001011000000101" => data <= "000000";
				when "001001011000000110" => data <= "000000";
				when "001001011000000111" => data <= "000000";
				when "001001011000001000" => data <= "000000";
				when "001001011000001001" => data <= "000000";
				when "001001011000001010" => data <= "000000";
				when "001001011000001011" => data <= "000000";
				when "001001011000001100" => data <= "000000";
				when "001001011000001101" => data <= "000000";
				when "001001011000001110" => data <= "000000";
				when "001001011000001111" => data <= "000000";
				when "001001011000010000" => data <= "000000";
				when "001001011000010001" => data <= "000000";
				when "001001011000010010" => data <= "000000";
				when "001001011000010011" => data <= "000000";
				when "001001011000010100" => data <= "000000";
				when "001001011000010101" => data <= "000000";
				when "001001011000010110" => data <= "000000";
				when "001001011000010111" => data <= "000000";
				when "001001011000011000" => data <= "000000";
				when "001001011000011001" => data <= "000000";
				when "001001011000011010" => data <= "000000";
				when "001001011000011011" => data <= "000000";
				when "001001011000011100" => data <= "000000";
				when "001001011000011101" => data <= "000000";
				when "001001011000011110" => data <= "000000";
				when "001001011000011111" => data <= "000000";
				when "001001011000100000" => data <= "000000";
				when "001001011000100001" => data <= "000000";
				when "001001011000100010" => data <= "000000";
				when "001001011000100011" => data <= "000000";
				when "001001011000100100" => data <= "000000";
				when "001001011000100101" => data <= "000000";
				when "001001011000100110" => data <= "000000";
				when "001001011000100111" => data <= "000000";
				when "001001011000101000" => data <= "000000";
				when "001001011000101001" => data <= "000000";
				when "001001011000101010" => data <= "000000";
				when "001001011000101011" => data <= "000000";
				when "001001011000101100" => data <= "000000";
				when "001001011000101101" => data <= "000000";
				when "001001011000101110" => data <= "000000";
				when "001001011000101111" => data <= "000000";
				when "001001011000110000" => data <= "000000";
				when "001001011000110001" => data <= "000000";
				when "001001011000110010" => data <= "000000";
				when "001001011000110011" => data <= "000000";
				when "001001011000110100" => data <= "000000";
				when "001001011000110101" => data <= "000000";
				when "001001011000110110" => data <= "000000";
				when "001001011000110111" => data <= "000000";
				when "001001011000111000" => data <= "000000";
				when "001001011000111001" => data <= "000000";
				when "001001011000111010" => data <= "000000";
				when "001001011000111011" => data <= "000000";
				when "001001011000111100" => data <= "000000";
				when "001001011000111101" => data <= "000000";
				when "001001011000111110" => data <= "000000";
				when "001001011000111111" => data <= "000000";
				when "001001011001000000" => data <= "000000";
				when "001001011001000001" => data <= "000000";
				when "001001011001000010" => data <= "000000";
				when "001001011001000011" => data <= "000000";
				when "001001011001000100" => data <= "000000";
				when "001001011001000101" => data <= "000000";
				when "001001011001000110" => data <= "000000";
				when "001001011001000111" => data <= "000000";
				when "001001011001001000" => data <= "000000";
				when "001001011001001001" => data <= "000000";
				when "001001011001001010" => data <= "000000";
				when "001001011001001011" => data <= "000000";
				when "001001011001001100" => data <= "000000";
				when "001001011001001101" => data <= "000000";
				when "001001011001001110" => data <= "000000";
				when "001001011001001111" => data <= "000000";
				when "001001011001010000" => data <= "000000";
				when "001001011001010001" => data <= "000000";
				when "001001011001010010" => data <= "000000";
				when "001001011001010011" => data <= "000000";
				when "001001011001010100" => data <= "000000";
				when "001001011001010101" => data <= "000000";
				when "001001011001010110" => data <= "000000";
				when "001001011001010111" => data <= "000000";
				when "001001011001011000" => data <= "000000";
				when "001001011001011001" => data <= "000000";
				when "001001011001011010" => data <= "000000";
				when "001001011001011011" => data <= "000000";
				when "001001011001011100" => data <= "000000";
				when "001001011001011101" => data <= "000000";
				when "001001011001011110" => data <= "000000";
				when "001001011001011111" => data <= "000000";
				when "001001011001100000" => data <= "000000";
				when "001001011001100001" => data <= "000000";
				when "001001011001100010" => data <= "000000";
				when "001001011001100011" => data <= "000000";
				when "001001011001100100" => data <= "000000";
				when "001001011001100101" => data <= "000000";
				when "001001011001100110" => data <= "000000";
				when "001001011001100111" => data <= "000000";
				when "001001011001101000" => data <= "000000";
				when "001001011001101001" => data <= "000000";
				when "001001011001101010" => data <= "000000";
				when "001001011001101011" => data <= "000000";
				when "001001011001101100" => data <= "000000";
				when "001001011001101101" => data <= "000000";
				when "001001011001101110" => data <= "000000";
				when "001001011001101111" => data <= "000000";
				when "001001011001110000" => data <= "000000";
				when "001001011001110001" => data <= "000000";
				when "001001011001110010" => data <= "000000";
				when "001001011001110011" => data <= "000000";
				when "001001011001110100" => data <= "000000";
				when "001001011001110101" => data <= "000000";
				when "001001011001110110" => data <= "000000";
				when "001001011001110111" => data <= "000000";
				when "001001011001111000" => data <= "000000";
				when "001001011001111001" => data <= "000000";
				when "001001011001111010" => data <= "000000";
				when "001001011001111011" => data <= "000000";
				when "001001011001111100" => data <= "000000";
				when "001001011001111101" => data <= "000000";
				when "001001011001111110" => data <= "000000";
				when "001001011001111111" => data <= "000000";
				when "001001011010000000" => data <= "000000";
				when "001001011010000001" => data <= "000000";
				when "001001011010000010" => data <= "000000";
				when "001001011010000011" => data <= "000000";
				when "001001011010000100" => data <= "000000";
				when "001001011010000101" => data <= "000000";
				when "001001011010000110" => data <= "000000";
				when "001001011010000111" => data <= "000000";
				when "001001011010001000" => data <= "000000";
				when "001001011010001001" => data <= "000000";
				when "001001011010001010" => data <= "000000";
				when "001001011010001011" => data <= "000000";
				when "001001011010001100" => data <= "000000";
				when "001001011010001101" => data <= "000000";
				when "001001011010001110" => data <= "000000";
				when "001001011010001111" => data <= "000000";
				when "001001011010010000" => data <= "000000";
				when "001001011010010001" => data <= "000000";
				when "001001011010010010" => data <= "000000";
				when "001001011010010011" => data <= "000000";
				when "001001011010010100" => data <= "000000";
				when "001001011010010101" => data <= "000000";
				when "001001011010010110" => data <= "000000";
				when "001001011010010111" => data <= "000000";
				when "001001011010011000" => data <= "000000";
				when "001001011010011001" => data <= "000000";
				when "001001011010011010" => data <= "000000";
				when "001001011010011011" => data <= "000000";
				when "001001011010011100" => data <= "000000";
				when "001001011010011101" => data <= "000000";
				when "001001011010011110" => data <= "000000";
				when "001001011010011111" => data <= "000000";
				when "001001100000000000" => data <= "000000";
				when "001001100000000001" => data <= "000000";
				when "001001100000000010" => data <= "000000";
				when "001001100000000011" => data <= "000000";
				when "001001100000000100" => data <= "000000";
				when "001001100000000101" => data <= "000000";
				when "001001100000000110" => data <= "000000";
				when "001001100000000111" => data <= "000000";
				when "001001100000001000" => data <= "000000";
				when "001001100000001001" => data <= "000000";
				when "001001100000001010" => data <= "000000";
				when "001001100000001011" => data <= "000000";
				when "001001100000001100" => data <= "000000";
				when "001001100000001101" => data <= "000000";
				when "001001100000001110" => data <= "000000";
				when "001001100000001111" => data <= "000000";
				when "001001100000010000" => data <= "000000";
				when "001001100000010001" => data <= "000000";
				when "001001100000010010" => data <= "000000";
				when "001001100000010011" => data <= "000000";
				when "001001100000010100" => data <= "000000";
				when "001001100000010101" => data <= "000000";
				when "001001100000010110" => data <= "000000";
				when "001001100000010111" => data <= "000000";
				when "001001100000011000" => data <= "000000";
				when "001001100000011001" => data <= "000000";
				when "001001100000011010" => data <= "000000";
				when "001001100000011011" => data <= "000000";
				when "001001100000011100" => data <= "000000";
				when "001001100000011101" => data <= "000000";
				when "001001100000011110" => data <= "000000";
				when "001001100000011111" => data <= "000000";
				when "001001100000100000" => data <= "000000";
				when "001001100000100001" => data <= "000000";
				when "001001100000100010" => data <= "000000";
				when "001001100000100011" => data <= "000000";
				when "001001100000100100" => data <= "000000";
				when "001001100000100101" => data <= "000000";
				when "001001100000100110" => data <= "000000";
				when "001001100000100111" => data <= "000000";
				when "001001100000101000" => data <= "000000";
				when "001001100000101001" => data <= "000000";
				when "001001100000101010" => data <= "000000";
				when "001001100000101011" => data <= "000000";
				when "001001100000101100" => data <= "000000";
				when "001001100000101101" => data <= "000000";
				when "001001100000101110" => data <= "000000";
				when "001001100000101111" => data <= "000000";
				when "001001100000110000" => data <= "000000";
				when "001001100000110001" => data <= "000000";
				when "001001100000110010" => data <= "000000";
				when "001001100000110011" => data <= "000000";
				when "001001100000110100" => data <= "000000";
				when "001001100000110101" => data <= "000000";
				when "001001100000110110" => data <= "000000";
				when "001001100000110111" => data <= "000000";
				when "001001100000111000" => data <= "000000";
				when "001001100000111001" => data <= "000000";
				when "001001100000111010" => data <= "000000";
				when "001001100000111011" => data <= "000000";
				when "001001100000111100" => data <= "000000";
				when "001001100000111101" => data <= "000000";
				when "001001100000111110" => data <= "000000";
				when "001001100000111111" => data <= "000000";
				when "001001100001000000" => data <= "000000";
				when "001001100001000001" => data <= "000000";
				when "001001100001000010" => data <= "000000";
				when "001001100001000011" => data <= "000000";
				when "001001100001000100" => data <= "000000";
				when "001001100001000101" => data <= "000000";
				when "001001100001000110" => data <= "000000";
				when "001001100001000111" => data <= "000000";
				when "001001100001001000" => data <= "000000";
				when "001001100001001001" => data <= "000000";
				when "001001100001001010" => data <= "000000";
				when "001001100001001011" => data <= "000000";
				when "001001100001001100" => data <= "000000";
				when "001001100001001101" => data <= "000000";
				when "001001100001001110" => data <= "000000";
				when "001001100001001111" => data <= "000000";
				when "001001100001010000" => data <= "000000";
				when "001001100001010001" => data <= "000000";
				when "001001100001010010" => data <= "000000";
				when "001001100001010011" => data <= "000000";
				when "001001100001010100" => data <= "000000";
				when "001001100001010101" => data <= "000000";
				when "001001100001010110" => data <= "000000";
				when "001001100001010111" => data <= "000000";
				when "001001100001011000" => data <= "000000";
				when "001001100001011001" => data <= "000000";
				when "001001100001011010" => data <= "000000";
				when "001001100001011011" => data <= "000000";
				when "001001100001011100" => data <= "000000";
				when "001001100001011101" => data <= "000000";
				when "001001100001011110" => data <= "000000";
				when "001001100001011111" => data <= "000000";
				when "001001100001100000" => data <= "000000";
				when "001001100001100001" => data <= "000000";
				when "001001100001100010" => data <= "000000";
				when "001001100001100011" => data <= "000000";
				when "001001100001100100" => data <= "000000";
				when "001001100001100101" => data <= "000000";
				when "001001100001100110" => data <= "000000";
				when "001001100001100111" => data <= "000000";
				when "001001100001101000" => data <= "000000";
				when "001001100001101001" => data <= "000000";
				when "001001100001101010" => data <= "000000";
				when "001001100001101011" => data <= "000000";
				when "001001100001101100" => data <= "000000";
				when "001001100001101101" => data <= "000000";
				when "001001100001101110" => data <= "000000";
				when "001001100001101111" => data <= "000000";
				when "001001100001110000" => data <= "000000";
				when "001001100001110001" => data <= "000000";
				when "001001100001110010" => data <= "000000";
				when "001001100001110011" => data <= "000000";
				when "001001100001110100" => data <= "000000";
				when "001001100001110101" => data <= "000000";
				when "001001100001110110" => data <= "000000";
				when "001001100001110111" => data <= "000000";
				when "001001100001111000" => data <= "000000";
				when "001001100001111001" => data <= "000000";
				when "001001100001111010" => data <= "000000";
				when "001001100001111011" => data <= "000000";
				when "001001100001111100" => data <= "000000";
				when "001001100001111101" => data <= "000000";
				when "001001100001111110" => data <= "000000";
				when "001001100001111111" => data <= "000000";
				when "001001100010000000" => data <= "000000";
				when "001001100010000001" => data <= "000000";
				when "001001100010000010" => data <= "000000";
				when "001001100010000011" => data <= "000000";
				when "001001100010000100" => data <= "000000";
				when "001001100010000101" => data <= "000000";
				when "001001100010000110" => data <= "000000";
				when "001001100010000111" => data <= "000000";
				when "001001100010001000" => data <= "000000";
				when "001001100010001001" => data <= "000000";
				when "001001100010001010" => data <= "000000";
				when "001001100010001011" => data <= "000000";
				when "001001100010001100" => data <= "000000";
				when "001001100010001101" => data <= "000000";
				when "001001100010001110" => data <= "000000";
				when "001001100010001111" => data <= "000000";
				when "001001100010010000" => data <= "000000";
				when "001001100010010001" => data <= "000000";
				when "001001100010010010" => data <= "000000";
				when "001001100010010011" => data <= "000000";
				when "001001100010010100" => data <= "000000";
				when "001001100010010101" => data <= "000000";
				when "001001100010010110" => data <= "000000";
				when "001001100010010111" => data <= "000000";
				when "001001100010011000" => data <= "000000";
				when "001001100010011001" => data <= "000000";
				when "001001100010011010" => data <= "000000";
				when "001001100010011011" => data <= "000000";
				when "001001100010011100" => data <= "000000";
				when "001001100010011101" => data <= "000000";
				when "001001100010011110" => data <= "000000";
				when "001001100010011111" => data <= "000000";
				when "001001101000000000" => data <= "000000";
				when "001001101000000001" => data <= "000000";
				when "001001101000000010" => data <= "000000";
				when "001001101000000011" => data <= "000000";
				when "001001101000000100" => data <= "000000";
				when "001001101000000101" => data <= "000000";
				when "001001101000000110" => data <= "000000";
				when "001001101000000111" => data <= "000000";
				when "001001101000001000" => data <= "000000";
				when "001001101000001001" => data <= "000000";
				when "001001101000001010" => data <= "000000";
				when "001001101000001011" => data <= "000000";
				when "001001101000001100" => data <= "000000";
				when "001001101000001101" => data <= "000000";
				when "001001101000001110" => data <= "000000";
				when "001001101000001111" => data <= "000000";
				when "001001101000010000" => data <= "000000";
				when "001001101000010001" => data <= "000000";
				when "001001101000010010" => data <= "000000";
				when "001001101000010011" => data <= "000000";
				when "001001101000010100" => data <= "000000";
				when "001001101000010101" => data <= "000000";
				when "001001101000010110" => data <= "000000";
				when "001001101000010111" => data <= "000000";
				when "001001101000011000" => data <= "000000";
				when "001001101000011001" => data <= "000000";
				when "001001101000011010" => data <= "000000";
				when "001001101000011011" => data <= "000000";
				when "001001101000011100" => data <= "000000";
				when "001001101000011101" => data <= "000000";
				when "001001101000011110" => data <= "000000";
				when "001001101000011111" => data <= "000000";
				when "001001101000100000" => data <= "000000";
				when "001001101000100001" => data <= "000000";
				when "001001101000100010" => data <= "000000";
				when "001001101000100011" => data <= "000000";
				when "001001101000100100" => data <= "000000";
				when "001001101000100101" => data <= "000000";
				when "001001101000100110" => data <= "000000";
				when "001001101000100111" => data <= "000000";
				when "001001101000101000" => data <= "000000";
				when "001001101000101001" => data <= "000000";
				when "001001101000101010" => data <= "000000";
				when "001001101000101011" => data <= "000000";
				when "001001101000101100" => data <= "000000";
				when "001001101000101101" => data <= "000000";
				when "001001101000101110" => data <= "000000";
				when "001001101000101111" => data <= "000000";
				when "001001101000110000" => data <= "000000";
				when "001001101000110001" => data <= "000000";
				when "001001101000110010" => data <= "000000";
				when "001001101000110011" => data <= "000000";
				when "001001101000110100" => data <= "000000";
				when "001001101000110101" => data <= "000000";
				when "001001101000110110" => data <= "000000";
				when "001001101000110111" => data <= "000000";
				when "001001101000111000" => data <= "000000";
				when "001001101000111001" => data <= "000000";
				when "001001101000111010" => data <= "000000";
				when "001001101000111011" => data <= "000000";
				when "001001101000111100" => data <= "000000";
				when "001001101000111101" => data <= "000000";
				when "001001101000111110" => data <= "000000";
				when "001001101000111111" => data <= "000000";
				when "001001101001000000" => data <= "000000";
				when "001001101001000001" => data <= "000000";
				when "001001101001000010" => data <= "000000";
				when "001001101001000011" => data <= "000000";
				when "001001101001000100" => data <= "000000";
				when "001001101001000101" => data <= "000000";
				when "001001101001000110" => data <= "000000";
				when "001001101001000111" => data <= "000000";
				when "001001101001001000" => data <= "000000";
				when "001001101001001001" => data <= "000000";
				when "001001101001001010" => data <= "000000";
				when "001001101001001011" => data <= "000000";
				when "001001101001001100" => data <= "000000";
				when "001001101001001101" => data <= "000000";
				when "001001101001001110" => data <= "000000";
				when "001001101001001111" => data <= "000000";
				when "001001101001010000" => data <= "000000";
				when "001001101001010001" => data <= "000000";
				when "001001101001010010" => data <= "000000";
				when "001001101001010011" => data <= "000000";
				when "001001101001010100" => data <= "000000";
				when "001001101001010101" => data <= "000000";
				when "001001101001010110" => data <= "000000";
				when "001001101001010111" => data <= "000000";
				when "001001101001011000" => data <= "000000";
				when "001001101001011001" => data <= "000000";
				when "001001101001011010" => data <= "000000";
				when "001001101001011011" => data <= "000000";
				when "001001101001011100" => data <= "000000";
				when "001001101001011101" => data <= "000000";
				when "001001101001011110" => data <= "000000";
				when "001001101001011111" => data <= "000000";
				when "001001101001100000" => data <= "000000";
				when "001001101001100001" => data <= "000000";
				when "001001101001100010" => data <= "000000";
				when "001001101001100011" => data <= "000000";
				when "001001101001100100" => data <= "000000";
				when "001001101001100101" => data <= "000000";
				when "001001101001100110" => data <= "000000";
				when "001001101001100111" => data <= "000000";
				when "001001101001101000" => data <= "000000";
				when "001001101001101001" => data <= "000000";
				when "001001101001101010" => data <= "000000";
				when "001001101001101011" => data <= "000000";
				when "001001101001101100" => data <= "000000";
				when "001001101001101101" => data <= "000000";
				when "001001101001101110" => data <= "000000";
				when "001001101001101111" => data <= "000000";
				when "001001101001110000" => data <= "000000";
				when "001001101001110001" => data <= "000000";
				when "001001101001110010" => data <= "000000";
				when "001001101001110011" => data <= "000000";
				when "001001101001110100" => data <= "000000";
				when "001001101001110101" => data <= "000000";
				when "001001101001110110" => data <= "000000";
				when "001001101001110111" => data <= "000000";
				when "001001101001111000" => data <= "000000";
				when "001001101001111001" => data <= "000000";
				when "001001101001111010" => data <= "000000";
				when "001001101001111011" => data <= "000000";
				when "001001101001111100" => data <= "000000";
				when "001001101001111101" => data <= "000000";
				when "001001101001111110" => data <= "000000";
				when "001001101001111111" => data <= "000000";
				when "001001101010000000" => data <= "000000";
				when "001001101010000001" => data <= "000000";
				when "001001101010000010" => data <= "000000";
				when "001001101010000011" => data <= "000000";
				when "001001101010000100" => data <= "000000";
				when "001001101010000101" => data <= "000000";
				when "001001101010000110" => data <= "000000";
				when "001001101010000111" => data <= "000000";
				when "001001101010001000" => data <= "000000";
				when "001001101010001001" => data <= "000000";
				when "001001101010001010" => data <= "000000";
				when "001001101010001011" => data <= "000000";
				when "001001101010001100" => data <= "000000";
				when "001001101010001101" => data <= "000000";
				when "001001101010001110" => data <= "000000";
				when "001001101010001111" => data <= "000000";
				when "001001101010010000" => data <= "000000";
				when "001001101010010001" => data <= "000000";
				when "001001101010010010" => data <= "000000";
				when "001001101010010011" => data <= "000000";
				when "001001101010010100" => data <= "000000";
				when "001001101010010101" => data <= "000000";
				when "001001101010010110" => data <= "000000";
				when "001001101010010111" => data <= "000000";
				when "001001101010011000" => data <= "000000";
				when "001001101010011001" => data <= "000000";
				when "001001101010011010" => data <= "000000";
				when "001001101010011011" => data <= "000000";
				when "001001101010011100" => data <= "000000";
				when "001001101010011101" => data <= "000000";
				when "001001101010011110" => data <= "000000";
				when "001001101010011111" => data <= "000000";
				when "001001110000000000" => data <= "000000";
				when "001001110000000001" => data <= "000000";
				when "001001110000000010" => data <= "000000";
				when "001001110000000011" => data <= "000000";
				when "001001110000000100" => data <= "000000";
				when "001001110000000101" => data <= "000000";
				when "001001110000000110" => data <= "000000";
				when "001001110000000111" => data <= "000000";
				when "001001110000001000" => data <= "000000";
				when "001001110000001001" => data <= "000000";
				when "001001110000001010" => data <= "000000";
				when "001001110000001011" => data <= "000000";
				when "001001110000001100" => data <= "000000";
				when "001001110000001101" => data <= "000000";
				when "001001110000001110" => data <= "000000";
				when "001001110000001111" => data <= "000000";
				when "001001110000010000" => data <= "000000";
				when "001001110000010001" => data <= "000000";
				when "001001110000010010" => data <= "000000";
				when "001001110000010011" => data <= "000000";
				when "001001110000010100" => data <= "000000";
				when "001001110000010101" => data <= "000000";
				when "001001110000010110" => data <= "000000";
				when "001001110000010111" => data <= "000000";
				when "001001110000011000" => data <= "000000";
				when "001001110000011001" => data <= "000000";
				when "001001110000011010" => data <= "000000";
				when "001001110000011011" => data <= "000000";
				when "001001110000011100" => data <= "000000";
				when "001001110000011101" => data <= "000000";
				when "001001110000011110" => data <= "000000";
				when "001001110000011111" => data <= "000000";
				when "001001110000100000" => data <= "000000";
				when "001001110000100001" => data <= "000000";
				when "001001110000100010" => data <= "000000";
				when "001001110000100011" => data <= "000000";
				when "001001110000100100" => data <= "000000";
				when "001001110000100101" => data <= "000000";
				when "001001110000100110" => data <= "000000";
				when "001001110000100111" => data <= "000000";
				when "001001110000101000" => data <= "000000";
				when "001001110000101001" => data <= "000000";
				when "001001110000101010" => data <= "000000";
				when "001001110000101011" => data <= "000000";
				when "001001110000101100" => data <= "000000";
				when "001001110000101101" => data <= "000000";
				when "001001110000101110" => data <= "000000";
				when "001001110000101111" => data <= "000000";
				when "001001110000110000" => data <= "000000";
				when "001001110000110001" => data <= "000000";
				when "001001110000110010" => data <= "000000";
				when "001001110000110011" => data <= "000000";
				when "001001110000110100" => data <= "000000";
				when "001001110000110101" => data <= "000000";
				when "001001110000110110" => data <= "000000";
				when "001001110000110111" => data <= "000000";
				when "001001110000111000" => data <= "000000";
				when "001001110000111001" => data <= "000000";
				when "001001110000111010" => data <= "000000";
				when "001001110000111011" => data <= "000000";
				when "001001110000111100" => data <= "000000";
				when "001001110000111101" => data <= "000000";
				when "001001110000111110" => data <= "000000";
				when "001001110000111111" => data <= "000000";
				when "001001110001000000" => data <= "000000";
				when "001001110001000001" => data <= "000000";
				when "001001110001000010" => data <= "000000";
				when "001001110001000011" => data <= "000000";
				when "001001110001000100" => data <= "000000";
				when "001001110001000101" => data <= "000000";
				when "001001110001000110" => data <= "000000";
				when "001001110001000111" => data <= "000000";
				when "001001110001001000" => data <= "000000";
				when "001001110001001001" => data <= "000000";
				when "001001110001001010" => data <= "000000";
				when "001001110001001011" => data <= "000000";
				when "001001110001001100" => data <= "000000";
				when "001001110001001101" => data <= "000000";
				when "001001110001001110" => data <= "000000";
				when "001001110001001111" => data <= "000000";
				when "001001110001010000" => data <= "000000";
				when "001001110001010001" => data <= "000000";
				when "001001110001010010" => data <= "000000";
				when "001001110001010011" => data <= "000000";
				when "001001110001010100" => data <= "000000";
				when "001001110001010101" => data <= "000000";
				when "001001110001010110" => data <= "000000";
				when "001001110001010111" => data <= "000000";
				when "001001110001011000" => data <= "000000";
				when "001001110001011001" => data <= "000000";
				when "001001110001011010" => data <= "000000";
				when "001001110001011011" => data <= "000000";
				when "001001110001011100" => data <= "000000";
				when "001001110001011101" => data <= "000000";
				when "001001110001011110" => data <= "000000";
				when "001001110001011111" => data <= "000000";
				when "001001110001100000" => data <= "000000";
				when "001001110001100001" => data <= "000000";
				when "001001110001100010" => data <= "000000";
				when "001001110001100011" => data <= "000000";
				when "001001110001100100" => data <= "000000";
				when "001001110001100101" => data <= "000000";
				when "001001110001100110" => data <= "000000";
				when "001001110001100111" => data <= "000000";
				when "001001110001101000" => data <= "000000";
				when "001001110001101001" => data <= "000000";
				when "001001110001101010" => data <= "000000";
				when "001001110001101011" => data <= "000000";
				when "001001110001101100" => data <= "000000";
				when "001001110001101101" => data <= "000000";
				when "001001110001101110" => data <= "000000";
				when "001001110001101111" => data <= "000000";
				when "001001110001110000" => data <= "000000";
				when "001001110001110001" => data <= "000000";
				when "001001110001110010" => data <= "000000";
				when "001001110001110011" => data <= "000000";
				when "001001110001110100" => data <= "000000";
				when "001001110001110101" => data <= "000000";
				when "001001110001110110" => data <= "000000";
				when "001001110001110111" => data <= "000000";
				when "001001110001111000" => data <= "000000";
				when "001001110001111001" => data <= "000000";
				when "001001110001111010" => data <= "000000";
				when "001001110001111011" => data <= "000000";
				when "001001110001111100" => data <= "000000";
				when "001001110001111101" => data <= "000000";
				when "001001110001111110" => data <= "000000";
				when "001001110001111111" => data <= "000000";
				when "001001110010000000" => data <= "000000";
				when "001001110010000001" => data <= "000000";
				when "001001110010000010" => data <= "000000";
				when "001001110010000011" => data <= "000000";
				when "001001110010000100" => data <= "000000";
				when "001001110010000101" => data <= "000000";
				when "001001110010000110" => data <= "000000";
				when "001001110010000111" => data <= "000000";
				when "001001110010001000" => data <= "000000";
				when "001001110010001001" => data <= "000000";
				when "001001110010001010" => data <= "000000";
				when "001001110010001011" => data <= "000000";
				when "001001110010001100" => data <= "000000";
				when "001001110010001101" => data <= "000000";
				when "001001110010001110" => data <= "000000";
				when "001001110010001111" => data <= "000000";
				when "001001110010010000" => data <= "000000";
				when "001001110010010001" => data <= "000000";
				when "001001110010010010" => data <= "000000";
				when "001001110010010011" => data <= "000000";
				when "001001110010010100" => data <= "000000";
				when "001001110010010101" => data <= "000000";
				when "001001110010010110" => data <= "000000";
				when "001001110010010111" => data <= "000000";
				when "001001110010011000" => data <= "000000";
				when "001001110010011001" => data <= "000000";
				when "001001110010011010" => data <= "000000";
				when "001001110010011011" => data <= "000000";
				when "001001110010011100" => data <= "000000";
				when "001001110010011101" => data <= "000000";
				when "001001110010011110" => data <= "000000";
				when "001001110010011111" => data <= "000000";
				when "001001111000000000" => data <= "000000";
				when "001001111000000001" => data <= "000000";
				when "001001111000000010" => data <= "000000";
				when "001001111000000011" => data <= "000000";
				when "001001111000000100" => data <= "000000";
				when "001001111000000101" => data <= "000000";
				when "001001111000000110" => data <= "000000";
				when "001001111000000111" => data <= "000000";
				when "001001111000001000" => data <= "000000";
				when "001001111000001001" => data <= "000000";
				when "001001111000001010" => data <= "000000";
				when "001001111000001011" => data <= "000000";
				when "001001111000001100" => data <= "000000";
				when "001001111000001101" => data <= "000000";
				when "001001111000001110" => data <= "000000";
				when "001001111000001111" => data <= "000000";
				when "001001111000010000" => data <= "000000";
				when "001001111000010001" => data <= "000000";
				when "001001111000010010" => data <= "000000";
				when "001001111000010011" => data <= "000000";
				when "001001111000010100" => data <= "000000";
				when "001001111000010101" => data <= "000000";
				when "001001111000010110" => data <= "000000";
				when "001001111000010111" => data <= "000000";
				when "001001111000011000" => data <= "000000";
				when "001001111000011001" => data <= "000000";
				when "001001111000011010" => data <= "000000";
				when "001001111000011011" => data <= "000000";
				when "001001111000011100" => data <= "000000";
				when "001001111000011101" => data <= "000000";
				when "001001111000011110" => data <= "000000";
				when "001001111000011111" => data <= "000000";
				when "001001111000100000" => data <= "000000";
				when "001001111000100001" => data <= "000000";
				when "001001111000100010" => data <= "000000";
				when "001001111000100011" => data <= "000000";
				when "001001111000100100" => data <= "000000";
				when "001001111000100101" => data <= "000000";
				when "001001111000100110" => data <= "000000";
				when "001001111000100111" => data <= "000000";
				when "001001111000101000" => data <= "000000";
				when "001001111000101001" => data <= "000000";
				when "001001111000101010" => data <= "000000";
				when "001001111000101011" => data <= "000000";
				when "001001111000101100" => data <= "000000";
				when "001001111000101101" => data <= "000000";
				when "001001111000101110" => data <= "000000";
				when "001001111000101111" => data <= "000000";
				when "001001111000110000" => data <= "000000";
				when "001001111000110001" => data <= "000000";
				when "001001111000110010" => data <= "000000";
				when "001001111000110011" => data <= "000000";
				when "001001111000110100" => data <= "000000";
				when "001001111000110101" => data <= "000000";
				when "001001111000110110" => data <= "000000";
				when "001001111000110111" => data <= "000000";
				when "001001111000111000" => data <= "000000";
				when "001001111000111001" => data <= "000000";
				when "001001111000111010" => data <= "000000";
				when "001001111000111011" => data <= "000000";
				when "001001111000111100" => data <= "000000";
				when "001001111000111101" => data <= "000000";
				when "001001111000111110" => data <= "000000";
				when "001001111000111111" => data <= "000000";
				when "001001111001000000" => data <= "000000";
				when "001001111001000001" => data <= "000000";
				when "001001111001000010" => data <= "000000";
				when "001001111001000011" => data <= "000000";
				when "001001111001000100" => data <= "000000";
				when "001001111001000101" => data <= "000000";
				when "001001111001000110" => data <= "000000";
				when "001001111001000111" => data <= "000000";
				when "001001111001001000" => data <= "000000";
				when "001001111001001001" => data <= "000000";
				when "001001111001001010" => data <= "000000";
				when "001001111001001011" => data <= "000000";
				when "001001111001001100" => data <= "000000";
				when "001001111001001101" => data <= "000000";
				when "001001111001001110" => data <= "000000";
				when "001001111001001111" => data <= "000000";
				when "001001111001010000" => data <= "000000";
				when "001001111001010001" => data <= "000000";
				when "001001111001010010" => data <= "000000";
				when "001001111001010011" => data <= "000000";
				when "001001111001010100" => data <= "000000";
				when "001001111001010101" => data <= "000000";
				when "001001111001010110" => data <= "000000";
				when "001001111001010111" => data <= "000000";
				when "001001111001011000" => data <= "000000";
				when "001001111001011001" => data <= "000000";
				when "001001111001011010" => data <= "000000";
				when "001001111001011011" => data <= "000000";
				when "001001111001011100" => data <= "000000";
				when "001001111001011101" => data <= "000000";
				when "001001111001011110" => data <= "000000";
				when "001001111001011111" => data <= "000000";
				when "001001111001100000" => data <= "000000";
				when "001001111001100001" => data <= "000000";
				when "001001111001100010" => data <= "000000";
				when "001001111001100011" => data <= "000000";
				when "001001111001100100" => data <= "000000";
				when "001001111001100101" => data <= "000000";
				when "001001111001100110" => data <= "000000";
				when "001001111001100111" => data <= "000000";
				when "001001111001101000" => data <= "000000";
				when "001001111001101001" => data <= "000000";
				when "001001111001101010" => data <= "000000";
				when "001001111001101011" => data <= "000000";
				when "001001111001101100" => data <= "000000";
				when "001001111001101101" => data <= "000000";
				when "001001111001101110" => data <= "000000";
				when "001001111001101111" => data <= "000000";
				when "001001111001110000" => data <= "000000";
				when "001001111001110001" => data <= "000000";
				when "001001111001110010" => data <= "000000";
				when "001001111001110011" => data <= "000000";
				when "001001111001110100" => data <= "000000";
				when "001001111001110101" => data <= "000000";
				when "001001111001110110" => data <= "000000";
				when "001001111001110111" => data <= "000000";
				when "001001111001111000" => data <= "000000";
				when "001001111001111001" => data <= "000000";
				when "001001111001111010" => data <= "000000";
				when "001001111001111011" => data <= "000000";
				when "001001111001111100" => data <= "000000";
				when "001001111001111101" => data <= "000000";
				when "001001111001111110" => data <= "000000";
				when "001001111001111111" => data <= "000000";
				when "001001111010000000" => data <= "000000";
				when "001001111010000001" => data <= "000000";
				when "001001111010000010" => data <= "000000";
				when "001001111010000011" => data <= "000000";
				when "001001111010000100" => data <= "000000";
				when "001001111010000101" => data <= "000000";
				when "001001111010000110" => data <= "000000";
				when "001001111010000111" => data <= "000000";
				when "001001111010001000" => data <= "000000";
				when "001001111010001001" => data <= "000000";
				when "001001111010001010" => data <= "000000";
				when "001001111010001011" => data <= "000000";
				when "001001111010001100" => data <= "000000";
				when "001001111010001101" => data <= "000000";
				when "001001111010001110" => data <= "000000";
				when "001001111010001111" => data <= "000000";
				when "001001111010010000" => data <= "000000";
				when "001001111010010001" => data <= "000000";
				when "001001111010010010" => data <= "000000";
				when "001001111010010011" => data <= "000000";
				when "001001111010010100" => data <= "000000";
				when "001001111010010101" => data <= "000000";
				when "001001111010010110" => data <= "000000";
				when "001001111010010111" => data <= "000000";
				when "001001111010011000" => data <= "000000";
				when "001001111010011001" => data <= "000000";
				when "001001111010011010" => data <= "000000";
				when "001001111010011011" => data <= "000000";
				when "001001111010011100" => data <= "000000";
				when "001001111010011101" => data <= "000000";
				when "001001111010011110" => data <= "000000";
				when "001001111010011111" => data <= "000000";
				when "001010000000000000" => data <= "000000";
				when "001010000000000001" => data <= "000000";
				when "001010000000000010" => data <= "000000";
				when "001010000000000011" => data <= "000000";
				when "001010000000000100" => data <= "000000";
				when "001010000000000101" => data <= "000000";
				when "001010000000000110" => data <= "000000";
				when "001010000000000111" => data <= "000000";
				when "001010000000001000" => data <= "000000";
				when "001010000000001001" => data <= "000000";
				when "001010000000001010" => data <= "000000";
				when "001010000000001011" => data <= "000000";
				when "001010000000001100" => data <= "000000";
				when "001010000000001101" => data <= "000000";
				when "001010000000001110" => data <= "000000";
				when "001010000000001111" => data <= "000000";
				when "001010000000010000" => data <= "000000";
				when "001010000000010001" => data <= "000000";
				when "001010000000010010" => data <= "000000";
				when "001010000000010011" => data <= "000000";
				when "001010000000010100" => data <= "000000";
				when "001010000000010101" => data <= "000000";
				when "001010000000010110" => data <= "000000";
				when "001010000000010111" => data <= "000000";
				when "001010000000011000" => data <= "000000";
				when "001010000000011001" => data <= "000000";
				when "001010000000011010" => data <= "000000";
				when "001010000000011011" => data <= "000000";
				when "001010000000011100" => data <= "000000";
				when "001010000000011101" => data <= "000000";
				when "001010000000011110" => data <= "000000";
				when "001010000000011111" => data <= "000000";
				when "001010000000100000" => data <= "000000";
				when "001010000000100001" => data <= "000000";
				when "001010000000100010" => data <= "000000";
				when "001010000000100011" => data <= "000000";
				when "001010000000100100" => data <= "000000";
				when "001010000000100101" => data <= "000000";
				when "001010000000100110" => data <= "000000";
				when "001010000000100111" => data <= "000000";
				when "001010000000101000" => data <= "000000";
				when "001010000000101001" => data <= "000000";
				when "001010000000101010" => data <= "000000";
				when "001010000000101011" => data <= "000000";
				when "001010000000101100" => data <= "000000";
				when "001010000000101101" => data <= "000000";
				when "001010000000101110" => data <= "000000";
				when "001010000000101111" => data <= "000000";
				when "001010000000110000" => data <= "000000";
				when "001010000000110001" => data <= "000000";
				when "001010000000110010" => data <= "000000";
				when "001010000000110011" => data <= "000000";
				when "001010000000110100" => data <= "000000";
				when "001010000000110101" => data <= "000000";
				when "001010000000110110" => data <= "000000";
				when "001010000000110111" => data <= "000000";
				when "001010000000111000" => data <= "000000";
				when "001010000000111001" => data <= "000000";
				when "001010000000111010" => data <= "000000";
				when "001010000000111011" => data <= "000000";
				when "001010000000111100" => data <= "000000";
				when "001010000000111101" => data <= "000000";
				when "001010000000111110" => data <= "000000";
				when "001010000000111111" => data <= "000000";
				when "001010000001000000" => data <= "000000";
				when "001010000001000001" => data <= "000000";
				when "001010000001000010" => data <= "000000";
				when "001010000001000011" => data <= "000000";
				when "001010000001000100" => data <= "000000";
				when "001010000001000101" => data <= "000000";
				when "001010000001000110" => data <= "000000";
				when "001010000001000111" => data <= "000000";
				when "001010000001001000" => data <= "000000";
				when "001010000001001001" => data <= "000000";
				when "001010000001001010" => data <= "000000";
				when "001010000001001011" => data <= "000000";
				when "001010000001001100" => data <= "000000";
				when "001010000001001101" => data <= "000000";
				when "001010000001001110" => data <= "000000";
				when "001010000001001111" => data <= "000000";
				when "001010000001010000" => data <= "000000";
				when "001010000001010001" => data <= "000000";
				when "001010000001010010" => data <= "000000";
				when "001010000001010011" => data <= "000000";
				when "001010000001010100" => data <= "000000";
				when "001010000001010101" => data <= "000000";
				when "001010000001010110" => data <= "000000";
				when "001010000001010111" => data <= "000000";
				when "001010000001011000" => data <= "000000";
				when "001010000001011001" => data <= "000000";
				when "001010000001011010" => data <= "000000";
				when "001010000001011011" => data <= "000000";
				when "001010000001011100" => data <= "000000";
				when "001010000001011101" => data <= "000000";
				when "001010000001011110" => data <= "000000";
				when "001010000001011111" => data <= "000000";
				when "001010000001100000" => data <= "000000";
				when "001010000001100001" => data <= "000000";
				when "001010000001100010" => data <= "000000";
				when "001010000001100011" => data <= "000000";
				when "001010000001100100" => data <= "000000";
				when "001010000001100101" => data <= "000000";
				when "001010000001100110" => data <= "000000";
				when "001010000001100111" => data <= "000000";
				when "001010000001101000" => data <= "000000";
				when "001010000001101001" => data <= "000000";
				when "001010000001101010" => data <= "000000";
				when "001010000001101011" => data <= "000000";
				when "001010000001101100" => data <= "000000";
				when "001010000001101101" => data <= "000000";
				when "001010000001101110" => data <= "000000";
				when "001010000001101111" => data <= "000000";
				when "001010000001110000" => data <= "000000";
				when "001010000001110001" => data <= "000000";
				when "001010000001110010" => data <= "000000";
				when "001010000001110011" => data <= "000000";
				when "001010000001110100" => data <= "000000";
				when "001010000001110101" => data <= "000000";
				when "001010000001110110" => data <= "000000";
				when "001010000001110111" => data <= "000000";
				when "001010000001111000" => data <= "000000";
				when "001010000001111001" => data <= "000000";
				when "001010000001111010" => data <= "000000";
				when "001010000001111011" => data <= "000000";
				when "001010000001111100" => data <= "000000";
				when "001010000001111101" => data <= "000000";
				when "001010000001111110" => data <= "000000";
				when "001010000001111111" => data <= "000000";
				when "001010000010000000" => data <= "000000";
				when "001010000010000001" => data <= "000000";
				when "001010000010000010" => data <= "000000";
				when "001010000010000011" => data <= "000000";
				when "001010000010000100" => data <= "000000";
				when "001010000010000101" => data <= "000000";
				when "001010000010000110" => data <= "000000";
				when "001010000010000111" => data <= "000000";
				when "001010000010001000" => data <= "000000";
				when "001010000010001001" => data <= "000000";
				when "001010000010001010" => data <= "000000";
				when "001010000010001011" => data <= "000000";
				when "001010000010001100" => data <= "000000";
				when "001010000010001101" => data <= "000000";
				when "001010000010001110" => data <= "000000";
				when "001010000010001111" => data <= "000000";
				when "001010000010010000" => data <= "000000";
				when "001010000010010001" => data <= "000000";
				when "001010000010010010" => data <= "000000";
				when "001010000010010011" => data <= "000000";
				when "001010000010010100" => data <= "000000";
				when "001010000010010101" => data <= "000000";
				when "001010000010010110" => data <= "000000";
				when "001010000010010111" => data <= "000000";
				when "001010000010011000" => data <= "000000";
				when "001010000010011001" => data <= "000000";
				when "001010000010011010" => data <= "000000";
				when "001010000010011011" => data <= "000000";
				when "001010000010011100" => data <= "000000";
				when "001010000010011101" => data <= "000000";
				when "001010000010011110" => data <= "000000";
				when "001010000010011111" => data <= "000000";
				when "001010001000000000" => data <= "000000";
				when "001010001000000001" => data <= "000000";
				when "001010001000000010" => data <= "000000";
				when "001010001000000011" => data <= "000000";
				when "001010001000000100" => data <= "000000";
				when "001010001000000101" => data <= "000000";
				when "001010001000000110" => data <= "000000";
				when "001010001000000111" => data <= "000000";
				when "001010001000001000" => data <= "000000";
				when "001010001000001001" => data <= "000000";
				when "001010001000001010" => data <= "000000";
				when "001010001000001011" => data <= "000000";
				when "001010001000001100" => data <= "000000";
				when "001010001000001101" => data <= "000000";
				when "001010001000001110" => data <= "000000";
				when "001010001000001111" => data <= "000000";
				when "001010001000010000" => data <= "000000";
				when "001010001000010001" => data <= "000000";
				when "001010001000010010" => data <= "000000";
				when "001010001000010011" => data <= "000000";
				when "001010001000010100" => data <= "000000";
				when "001010001000010101" => data <= "000000";
				when "001010001000010110" => data <= "000000";
				when "001010001000010111" => data <= "000000";
				when "001010001000011000" => data <= "000000";
				when "001010001000011001" => data <= "000000";
				when "001010001000011010" => data <= "000000";
				when "001010001000011011" => data <= "000000";
				when "001010001000011100" => data <= "000000";
				when "001010001000011101" => data <= "000000";
				when "001010001000011110" => data <= "000000";
				when "001010001000011111" => data <= "000000";
				when "001010001000100000" => data <= "000000";
				when "001010001000100001" => data <= "000000";
				when "001010001000100010" => data <= "000000";
				when "001010001000100011" => data <= "000000";
				when "001010001000100100" => data <= "000000";
				when "001010001000100101" => data <= "000000";
				when "001010001000100110" => data <= "000000";
				when "001010001000100111" => data <= "000000";
				when "001010001000101000" => data <= "000000";
				when "001010001000101001" => data <= "000000";
				when "001010001000101010" => data <= "000000";
				when "001010001000101011" => data <= "000000";
				when "001010001000101100" => data <= "000000";
				when "001010001000101101" => data <= "000000";
				when "001010001000101110" => data <= "000000";
				when "001010001000101111" => data <= "000000";
				when "001010001000110000" => data <= "000000";
				when "001010001000110001" => data <= "000000";
				when "001010001000110010" => data <= "000000";
				when "001010001000110011" => data <= "000000";
				when "001010001000110100" => data <= "000000";
				when "001010001000110101" => data <= "000000";
				when "001010001000110110" => data <= "000000";
				when "001010001000110111" => data <= "000000";
				when "001010001000111000" => data <= "000000";
				when "001010001000111001" => data <= "000000";
				when "001010001000111010" => data <= "000000";
				when "001010001000111011" => data <= "000000";
				when "001010001000111100" => data <= "000000";
				when "001010001000111101" => data <= "000000";
				when "001010001000111110" => data <= "000000";
				when "001010001000111111" => data <= "000000";
				when "001010001001000000" => data <= "000000";
				when "001010001001000001" => data <= "000000";
				when "001010001001000010" => data <= "000000";
				when "001010001001000011" => data <= "000000";
				when "001010001001000100" => data <= "000000";
				when "001010001001000101" => data <= "000000";
				when "001010001001000110" => data <= "000000";
				when "001010001001000111" => data <= "000000";
				when "001010001001001000" => data <= "000000";
				when "001010001001001001" => data <= "000000";
				when "001010001001001010" => data <= "000000";
				when "001010001001001011" => data <= "000000";
				when "001010001001001100" => data <= "000000";
				when "001010001001001101" => data <= "000000";
				when "001010001001001110" => data <= "000000";
				when "001010001001001111" => data <= "000000";
				when "001010001001010000" => data <= "000000";
				when "001010001001010001" => data <= "000000";
				when "001010001001010010" => data <= "000000";
				when "001010001001010011" => data <= "000000";
				when "001010001001010100" => data <= "000000";
				when "001010001001010101" => data <= "000000";
				when "001010001001010110" => data <= "000000";
				when "001010001001010111" => data <= "000000";
				when "001010001001011000" => data <= "000000";
				when "001010001001011001" => data <= "000000";
				when "001010001001011010" => data <= "000000";
				when "001010001001011011" => data <= "000000";
				when "001010001001011100" => data <= "000000";
				when "001010001001011101" => data <= "000000";
				when "001010001001011110" => data <= "000000";
				when "001010001001011111" => data <= "000000";
				when "001010001001100000" => data <= "000000";
				when "001010001001100001" => data <= "000000";
				when "001010001001100010" => data <= "000000";
				when "001010001001100011" => data <= "000000";
				when "001010001001100100" => data <= "000000";
				when "001010001001100101" => data <= "000000";
				when "001010001001100110" => data <= "000000";
				when "001010001001100111" => data <= "000000";
				when "001010001001101000" => data <= "000000";
				when "001010001001101001" => data <= "000000";
				when "001010001001101010" => data <= "000000";
				when "001010001001101011" => data <= "000000";
				when "001010001001101100" => data <= "000000";
				when "001010001001101101" => data <= "000000";
				when "001010001001101110" => data <= "000000";
				when "001010001001101111" => data <= "000000";
				when "001010001001110000" => data <= "000000";
				when "001010001001110001" => data <= "000000";
				when "001010001001110010" => data <= "000000";
				when "001010001001110011" => data <= "000000";
				when "001010001001110100" => data <= "000000";
				when "001010001001110101" => data <= "000000";
				when "001010001001110110" => data <= "000000";
				when "001010001001110111" => data <= "000000";
				when "001010001001111000" => data <= "000000";
				when "001010001001111001" => data <= "000000";
				when "001010001001111010" => data <= "000000";
				when "001010001001111011" => data <= "000000";
				when "001010001001111100" => data <= "000000";
				when "001010001001111101" => data <= "000000";
				when "001010001001111110" => data <= "000000";
				when "001010001001111111" => data <= "000000";
				when "001010001010000000" => data <= "000000";
				when "001010001010000001" => data <= "000000";
				when "001010001010000010" => data <= "000000";
				when "001010001010000011" => data <= "000000";
				when "001010001010000100" => data <= "000000";
				when "001010001010000101" => data <= "000000";
				when "001010001010000110" => data <= "000000";
				when "001010001010000111" => data <= "000000";
				when "001010001010001000" => data <= "000000";
				when "001010001010001001" => data <= "000000";
				when "001010001010001010" => data <= "000000";
				when "001010001010001011" => data <= "000000";
				when "001010001010001100" => data <= "000000";
				when "001010001010001101" => data <= "000000";
				when "001010001010001110" => data <= "000000";
				when "001010001010001111" => data <= "000000";
				when "001010001010010000" => data <= "000000";
				when "001010001010010001" => data <= "000000";
				when "001010001010010010" => data <= "000000";
				when "001010001010010011" => data <= "000000";
				when "001010001010010100" => data <= "000000";
				when "001010001010010101" => data <= "000000";
				when "001010001010010110" => data <= "000000";
				when "001010001010010111" => data <= "000000";
				when "001010001010011000" => data <= "000000";
				when "001010001010011001" => data <= "000000";
				when "001010001010011010" => data <= "000000";
				when "001010001010011011" => data <= "000000";
				when "001010001010011100" => data <= "000000";
				when "001010001010011101" => data <= "000000";
				when "001010001010011110" => data <= "000000";
				when "001010001010011111" => data <= "000000";
				when "001010010000000000" => data <= "000000";
				when "001010010000000001" => data <= "000000";
				when "001010010000000010" => data <= "000000";
				when "001010010000000011" => data <= "000000";
				when "001010010000000100" => data <= "000000";
				when "001010010000000101" => data <= "000000";
				when "001010010000000110" => data <= "000000";
				when "001010010000000111" => data <= "000000";
				when "001010010000001000" => data <= "000000";
				when "001010010000001001" => data <= "000000";
				when "001010010000001010" => data <= "000000";
				when "001010010000001011" => data <= "000000";
				when "001010010000001100" => data <= "000000";
				when "001010010000001101" => data <= "000000";
				when "001010010000001110" => data <= "000000";
				when "001010010000001111" => data <= "000000";
				when "001010010000010000" => data <= "000000";
				when "001010010000010001" => data <= "000000";
				when "001010010000010010" => data <= "000000";
				when "001010010000010011" => data <= "000000";
				when "001010010000010100" => data <= "000000";
				when "001010010000010101" => data <= "000000";
				when "001010010000010110" => data <= "000000";
				when "001010010000010111" => data <= "000000";
				when "001010010000011000" => data <= "000000";
				when "001010010000011001" => data <= "000000";
				when "001010010000011010" => data <= "000000";
				when "001010010000011011" => data <= "000000";
				when "001010010000011100" => data <= "000000";
				when "001010010000011101" => data <= "000000";
				when "001010010000011110" => data <= "000000";
				when "001010010000011111" => data <= "000000";
				when "001010010000100000" => data <= "000000";
				when "001010010000100001" => data <= "000000";
				when "001010010000100010" => data <= "000000";
				when "001010010000100011" => data <= "000000";
				when "001010010000100100" => data <= "000000";
				when "001010010000100101" => data <= "000000";
				when "001010010000100110" => data <= "000000";
				when "001010010000100111" => data <= "000000";
				when "001010010000101000" => data <= "000000";
				when "001010010000101001" => data <= "000000";
				when "001010010000101010" => data <= "000000";
				when "001010010000101011" => data <= "000000";
				when "001010010000101100" => data <= "000000";
				when "001010010000101101" => data <= "000000";
				when "001010010000101110" => data <= "000000";
				when "001010010000101111" => data <= "000000";
				when "001010010000110000" => data <= "000000";
				when "001010010000110001" => data <= "000000";
				when "001010010000110010" => data <= "000000";
				when "001010010000110011" => data <= "000000";
				when "001010010000110100" => data <= "000000";
				when "001010010000110101" => data <= "000000";
				when "001010010000110110" => data <= "000000";
				when "001010010000110111" => data <= "000000";
				when "001010010000111000" => data <= "000000";
				when "001010010000111001" => data <= "000000";
				when "001010010000111010" => data <= "000000";
				when "001010010000111011" => data <= "000000";
				when "001010010000111100" => data <= "000000";
				when "001010010000111101" => data <= "000000";
				when "001010010000111110" => data <= "000000";
				when "001010010000111111" => data <= "000000";
				when "001010010001000000" => data <= "000000";
				when "001010010001000001" => data <= "000000";
				when "001010010001000010" => data <= "000000";
				when "001010010001000011" => data <= "000000";
				when "001010010001000100" => data <= "000000";
				when "001010010001000101" => data <= "000000";
				when "001010010001000110" => data <= "000000";
				when "001010010001000111" => data <= "000000";
				when "001010010001001000" => data <= "000000";
				when "001010010001001001" => data <= "000000";
				when "001010010001001010" => data <= "000000";
				when "001010010001001011" => data <= "000000";
				when "001010010001001100" => data <= "000000";
				when "001010010001001101" => data <= "000000";
				when "001010010001001110" => data <= "000000";
				when "001010010001001111" => data <= "000000";
				when "001010010001010000" => data <= "000000";
				when "001010010001010001" => data <= "000000";
				when "001010010001010010" => data <= "000000";
				when "001010010001010011" => data <= "000000";
				when "001010010001010100" => data <= "000000";
				when "001010010001010101" => data <= "000000";
				when "001010010001010110" => data <= "000000";
				when "001010010001010111" => data <= "000000";
				when "001010010001011000" => data <= "000000";
				when "001010010001011001" => data <= "000000";
				when "001010010001011010" => data <= "000000";
				when "001010010001011011" => data <= "000000";
				when "001010010001011100" => data <= "000000";
				when "001010010001011101" => data <= "000000";
				when "001010010001011110" => data <= "000000";
				when "001010010001011111" => data <= "000000";
				when "001010010001100000" => data <= "000000";
				when "001010010001100001" => data <= "000000";
				when "001010010001100010" => data <= "000000";
				when "001010010001100011" => data <= "000000";
				when "001010010001100100" => data <= "000000";
				when "001010010001100101" => data <= "000000";
				when "001010010001100110" => data <= "000000";
				when "001010010001100111" => data <= "000000";
				when "001010010001101000" => data <= "000000";
				when "001010010001101001" => data <= "000000";
				when "001010010001101010" => data <= "000000";
				when "001010010001101011" => data <= "000000";
				when "001010010001101100" => data <= "000000";
				when "001010010001101101" => data <= "000000";
				when "001010010001101110" => data <= "000000";
				when "001010010001101111" => data <= "000000";
				when "001010010001110000" => data <= "000000";
				when "001010010001110001" => data <= "000000";
				when "001010010001110010" => data <= "000000";
				when "001010010001110011" => data <= "000000";
				when "001010010001110100" => data <= "000000";
				when "001010010001110101" => data <= "000000";
				when "001010010001110110" => data <= "000000";
				when "001010010001110111" => data <= "000000";
				when "001010010001111000" => data <= "000000";
				when "001010010001111001" => data <= "000000";
				when "001010010001111010" => data <= "000000";
				when "001010010001111011" => data <= "000000";
				when "001010010001111100" => data <= "000000";
				when "001010010001111101" => data <= "000000";
				when "001010010001111110" => data <= "000000";
				when "001010010001111111" => data <= "000000";
				when "001010010010000000" => data <= "000000";
				when "001010010010000001" => data <= "000000";
				when "001010010010000010" => data <= "000000";
				when "001010010010000011" => data <= "000000";
				when "001010010010000100" => data <= "000000";
				when "001010010010000101" => data <= "000000";
				when "001010010010000110" => data <= "000000";
				when "001010010010000111" => data <= "000000";
				when "001010010010001000" => data <= "000000";
				when "001010010010001001" => data <= "000000";
				when "001010010010001010" => data <= "000000";
				when "001010010010001011" => data <= "000000";
				when "001010010010001100" => data <= "000000";
				when "001010010010001101" => data <= "000000";
				when "001010010010001110" => data <= "000000";
				when "001010010010001111" => data <= "000000";
				when "001010010010010000" => data <= "000000";
				when "001010010010010001" => data <= "000000";
				when "001010010010010010" => data <= "000000";
				when "001010010010010011" => data <= "000000";
				when "001010010010010100" => data <= "000000";
				when "001010010010010101" => data <= "000000";
				when "001010010010010110" => data <= "000000";
				when "001010010010010111" => data <= "000000";
				when "001010010010011000" => data <= "000000";
				when "001010010010011001" => data <= "000000";
				when "001010010010011010" => data <= "000000";
				when "001010010010011011" => data <= "000000";
				when "001010010010011100" => data <= "000000";
				when "001010010010011101" => data <= "000000";
				when "001010010010011110" => data <= "000000";
				when "001010010010011111" => data <= "000000";
				when "001010011000000000" => data <= "000000";
				when "001010011000000001" => data <= "000000";
				when "001010011000000010" => data <= "000000";
				when "001010011000000011" => data <= "000000";
				when "001010011000000100" => data <= "000000";
				when "001010011000000101" => data <= "000000";
				when "001010011000000110" => data <= "000000";
				when "001010011000000111" => data <= "000000";
				when "001010011000001000" => data <= "000000";
				when "001010011000001001" => data <= "000000";
				when "001010011000001010" => data <= "000000";
				when "001010011000001011" => data <= "000000";
				when "001010011000001100" => data <= "000000";
				when "001010011000001101" => data <= "000000";
				when "001010011000001110" => data <= "000000";
				when "001010011000001111" => data <= "000000";
				when "001010011000010000" => data <= "000000";
				when "001010011000010001" => data <= "000000";
				when "001010011000010010" => data <= "000000";
				when "001010011000010011" => data <= "000000";
				when "001010011000010100" => data <= "000000";
				when "001010011000010101" => data <= "000000";
				when "001010011000010110" => data <= "000000";
				when "001010011000010111" => data <= "000000";
				when "001010011000011000" => data <= "000000";
				when "001010011000011001" => data <= "000000";
				when "001010011000011010" => data <= "000000";
				when "001010011000011011" => data <= "000000";
				when "001010011000011100" => data <= "000000";
				when "001010011000011101" => data <= "000000";
				when "001010011000011110" => data <= "000000";
				when "001010011000011111" => data <= "000000";
				when "001010011000100000" => data <= "000000";
				when "001010011000100001" => data <= "000000";
				when "001010011000100010" => data <= "000000";
				when "001010011000100011" => data <= "000000";
				when "001010011000100100" => data <= "000000";
				when "001010011000100101" => data <= "000000";
				when "001010011000100110" => data <= "000000";
				when "001010011000100111" => data <= "000000";
				when "001010011000101000" => data <= "000000";
				when "001010011000101001" => data <= "000000";
				when "001010011000101010" => data <= "000000";
				when "001010011000101011" => data <= "000000";
				when "001010011000101100" => data <= "000000";
				when "001010011000101101" => data <= "000000";
				when "001010011000101110" => data <= "000000";
				when "001010011000101111" => data <= "000000";
				when "001010011000110000" => data <= "000000";
				when "001010011000110001" => data <= "000000";
				when "001010011000110010" => data <= "000000";
				when "001010011000110011" => data <= "000000";
				when "001010011000110100" => data <= "000000";
				when "001010011000110101" => data <= "000000";
				when "001010011000110110" => data <= "000000";
				when "001010011000110111" => data <= "000000";
				when "001010011000111000" => data <= "000000";
				when "001010011000111001" => data <= "000000";
				when "001010011000111010" => data <= "000000";
				when "001010011000111011" => data <= "000000";
				when "001010011000111100" => data <= "000000";
				when "001010011000111101" => data <= "000000";
				when "001010011000111110" => data <= "000000";
				when "001010011000111111" => data <= "000000";
				when "001010011001000000" => data <= "000000";
				when "001010011001000001" => data <= "000000";
				when "001010011001000010" => data <= "000000";
				when "001010011001000011" => data <= "000000";
				when "001010011001000100" => data <= "000000";
				when "001010011001000101" => data <= "000000";
				when "001010011001000110" => data <= "000000";
				when "001010011001000111" => data <= "000000";
				when "001010011001001000" => data <= "000000";
				when "001010011001001001" => data <= "000000";
				when "001010011001001010" => data <= "000000";
				when "001010011001001011" => data <= "000000";
				when "001010011001001100" => data <= "000000";
				when "001010011001001101" => data <= "000000";
				when "001010011001001110" => data <= "000000";
				when "001010011001001111" => data <= "000000";
				when "001010011001010000" => data <= "000000";
				when "001010011001010001" => data <= "000000";
				when "001010011001010010" => data <= "000000";
				when "001010011001010011" => data <= "000000";
				when "001010011001010100" => data <= "000000";
				when "001010011001010101" => data <= "000000";
				when "001010011001010110" => data <= "000000";
				when "001010011001010111" => data <= "000000";
				when "001010011001011000" => data <= "000000";
				when "001010011001011001" => data <= "000000";
				when "001010011001011010" => data <= "000000";
				when "001010011001011011" => data <= "000000";
				when "001010011001011100" => data <= "000000";
				when "001010011001011101" => data <= "000000";
				when "001010011001011110" => data <= "000000";
				when "001010011001011111" => data <= "000000";
				when "001010011001100000" => data <= "000000";
				when "001010011001100001" => data <= "000000";
				when "001010011001100010" => data <= "000000";
				when "001010011001100011" => data <= "000000";
				when "001010011001100100" => data <= "000000";
				when "001010011001100101" => data <= "000000";
				when "001010011001100110" => data <= "000000";
				when "001010011001100111" => data <= "000000";
				when "001010011001101000" => data <= "000000";
				when "001010011001101001" => data <= "000000";
				when "001010011001101010" => data <= "000000";
				when "001010011001101011" => data <= "000000";
				when "001010011001101100" => data <= "000000";
				when "001010011001101101" => data <= "000000";
				when "001010011001101110" => data <= "000000";
				when "001010011001101111" => data <= "000000";
				when "001010011001110000" => data <= "000000";
				when "001010011001110001" => data <= "000000";
				when "001010011001110010" => data <= "000000";
				when "001010011001110011" => data <= "000000";
				when "001010011001110100" => data <= "000000";
				when "001010011001110101" => data <= "000000";
				when "001010011001110110" => data <= "000000";
				when "001010011001110111" => data <= "000000";
				when "001010011001111000" => data <= "000000";
				when "001010011001111001" => data <= "000000";
				when "001010011001111010" => data <= "000000";
				when "001010011001111011" => data <= "000000";
				when "001010011001111100" => data <= "000000";
				when "001010011001111101" => data <= "000000";
				when "001010011001111110" => data <= "000000";
				when "001010011001111111" => data <= "000000";
				when "001010011010000000" => data <= "000000";
				when "001010011010000001" => data <= "000000";
				when "001010011010000010" => data <= "000000";
				when "001010011010000011" => data <= "000000";
				when "001010011010000100" => data <= "000000";
				when "001010011010000101" => data <= "000000";
				when "001010011010000110" => data <= "000000";
				when "001010011010000111" => data <= "000000";
				when "001010011010001000" => data <= "000000";
				when "001010011010001001" => data <= "000000";
				when "001010011010001010" => data <= "000000";
				when "001010011010001011" => data <= "000000";
				when "001010011010001100" => data <= "000000";
				when "001010011010001101" => data <= "000000";
				when "001010011010001110" => data <= "000000";
				when "001010011010001111" => data <= "000000";
				when "001010011010010000" => data <= "000000";
				when "001010011010010001" => data <= "000000";
				when "001010011010010010" => data <= "000000";
				when "001010011010010011" => data <= "000000";
				when "001010011010010100" => data <= "000000";
				when "001010011010010101" => data <= "000000";
				when "001010011010010110" => data <= "000000";
				when "001010011010010111" => data <= "000000";
				when "001010011010011000" => data <= "000000";
				when "001010011010011001" => data <= "000000";
				when "001010011010011010" => data <= "000000";
				when "001010011010011011" => data <= "000000";
				when "001010011010011100" => data <= "000000";
				when "001010011010011101" => data <= "000000";
				when "001010011010011110" => data <= "000000";
				when "001010011010011111" => data <= "000000";
				when "001010100000000000" => data <= "000000";
				when "001010100000000001" => data <= "000000";
				when "001010100000000010" => data <= "000000";
				when "001010100000000011" => data <= "000000";
				when "001010100000000100" => data <= "000000";
				when "001010100000000101" => data <= "000000";
				when "001010100000000110" => data <= "000000";
				when "001010100000000111" => data <= "000000";
				when "001010100000001000" => data <= "000000";
				when "001010100000001001" => data <= "000000";
				when "001010100000001010" => data <= "000000";
				when "001010100000001011" => data <= "000000";
				when "001010100000001100" => data <= "000000";
				when "001010100000001101" => data <= "000000";
				when "001010100000001110" => data <= "000000";
				when "001010100000001111" => data <= "000000";
				when "001010100000010000" => data <= "000000";
				when "001010100000010001" => data <= "000000";
				when "001010100000010010" => data <= "000000";
				when "001010100000010011" => data <= "000000";
				when "001010100000010100" => data <= "000000";
				when "001010100000010101" => data <= "000000";
				when "001010100000010110" => data <= "000000";
				when "001010100000010111" => data <= "000000";
				when "001010100000011000" => data <= "000000";
				when "001010100000011001" => data <= "000000";
				when "001010100000011010" => data <= "000000";
				when "001010100000011011" => data <= "000000";
				when "001010100000011100" => data <= "000000";
				when "001010100000011101" => data <= "000000";
				when "001010100000011110" => data <= "000000";
				when "001010100000011111" => data <= "000000";
				when "001010100000100000" => data <= "000000";
				when "001010100000100001" => data <= "000000";
				when "001010100000100010" => data <= "000000";
				when "001010100000100011" => data <= "000000";
				when "001010100000100100" => data <= "000000";
				when "001010100000100101" => data <= "000000";
				when "001010100000100110" => data <= "000000";
				when "001010100000100111" => data <= "000000";
				when "001010100000101000" => data <= "000000";
				when "001010100000101001" => data <= "000000";
				when "001010100000101010" => data <= "000000";
				when "001010100000101011" => data <= "000000";
				when "001010100000101100" => data <= "000000";
				when "001010100000101101" => data <= "000000";
				when "001010100000101110" => data <= "000000";
				when "001010100000101111" => data <= "000000";
				when "001010100000110000" => data <= "000000";
				when "001010100000110001" => data <= "000000";
				when "001010100000110010" => data <= "000000";
				when "001010100000110011" => data <= "000000";
				when "001010100000110100" => data <= "000000";
				when "001010100000110101" => data <= "000000";
				when "001010100000110110" => data <= "000000";
				when "001010100000110111" => data <= "000000";
				when "001010100000111000" => data <= "000000";
				when "001010100000111001" => data <= "000000";
				when "001010100000111010" => data <= "000000";
				when "001010100000111011" => data <= "000000";
				when "001010100000111100" => data <= "000000";
				when "001010100000111101" => data <= "000000";
				when "001010100000111110" => data <= "000000";
				when "001010100000111111" => data <= "000000";
				when "001010100001000000" => data <= "000000";
				when "001010100001000001" => data <= "000000";
				when "001010100001000010" => data <= "000000";
				when "001010100001000011" => data <= "000000";
				when "001010100001000100" => data <= "000000";
				when "001010100001000101" => data <= "000000";
				when "001010100001000110" => data <= "000000";
				when "001010100001000111" => data <= "000000";
				when "001010100001001000" => data <= "000000";
				when "001010100001001001" => data <= "000000";
				when "001010100001001010" => data <= "000000";
				when "001010100001001011" => data <= "000000";
				when "001010100001001100" => data <= "000000";
				when "001010100001001101" => data <= "000000";
				when "001010100001001110" => data <= "000000";
				when "001010100001001111" => data <= "000000";
				when "001010100001010000" => data <= "000000";
				when "001010100001010001" => data <= "000000";
				when "001010100001010010" => data <= "000000";
				when "001010100001010011" => data <= "000000";
				when "001010100001010100" => data <= "000000";
				when "001010100001010101" => data <= "000000";
				when "001010100001010110" => data <= "000000";
				when "001010100001010111" => data <= "000000";
				when "001010100001011000" => data <= "000000";
				when "001010100001011001" => data <= "000000";
				when "001010100001011010" => data <= "000000";
				when "001010100001011011" => data <= "000000";
				when "001010100001011100" => data <= "000000";
				when "001010100001011101" => data <= "000000";
				when "001010100001011110" => data <= "000000";
				when "001010100001011111" => data <= "000000";
				when "001010100001100000" => data <= "000000";
				when "001010100001100001" => data <= "000000";
				when "001010100001100010" => data <= "000000";
				when "001010100001100011" => data <= "000000";
				when "001010100001100100" => data <= "000000";
				when "001010100001100101" => data <= "000000";
				when "001010100001100110" => data <= "000000";
				when "001010100001100111" => data <= "000000";
				when "001010100001101000" => data <= "000000";
				when "001010100001101001" => data <= "000000";
				when "001010100001101010" => data <= "000000";
				when "001010100001101011" => data <= "000000";
				when "001010100001101100" => data <= "000000";
				when "001010100001101101" => data <= "000000";
				when "001010100001101110" => data <= "000000";
				when "001010100001101111" => data <= "000000";
				when "001010100001110000" => data <= "000000";
				when "001010100001110001" => data <= "000000";
				when "001010100001110010" => data <= "000000";
				when "001010100001110011" => data <= "000000";
				when "001010100001110100" => data <= "000000";
				when "001010100001110101" => data <= "000000";
				when "001010100001110110" => data <= "000000";
				when "001010100001110111" => data <= "000000";
				when "001010100001111000" => data <= "000000";
				when "001010100001111001" => data <= "000000";
				when "001010100001111010" => data <= "000000";
				when "001010100001111011" => data <= "000000";
				when "001010100001111100" => data <= "000000";
				when "001010100001111101" => data <= "000000";
				when "001010100001111110" => data <= "000000";
				when "001010100001111111" => data <= "000000";
				when "001010100010000000" => data <= "000000";
				when "001010100010000001" => data <= "000000";
				when "001010100010000010" => data <= "000000";
				when "001010100010000011" => data <= "000000";
				when "001010100010000100" => data <= "000000";
				when "001010100010000101" => data <= "000000";
				when "001010100010000110" => data <= "000000";
				when "001010100010000111" => data <= "000000";
				when "001010100010001000" => data <= "000000";
				when "001010100010001001" => data <= "000000";
				when "001010100010001010" => data <= "000000";
				when "001010100010001011" => data <= "000000";
				when "001010100010001100" => data <= "000000";
				when "001010100010001101" => data <= "000000";
				when "001010100010001110" => data <= "000000";
				when "001010100010001111" => data <= "000000";
				when "001010100010010000" => data <= "000000";
				when "001010100010010001" => data <= "000000";
				when "001010100010010010" => data <= "000000";
				when "001010100010010011" => data <= "000000";
				when "001010100010010100" => data <= "000000";
				when "001010100010010101" => data <= "000000";
				when "001010100010010110" => data <= "000000";
				when "001010100010010111" => data <= "000000";
				when "001010100010011000" => data <= "000000";
				when "001010100010011001" => data <= "000000";
				when "001010100010011010" => data <= "000000";
				when "001010100010011011" => data <= "000000";
				when "001010100010011100" => data <= "000000";
				when "001010100010011101" => data <= "000000";
				when "001010100010011110" => data <= "000000";
				when "001010100010011111" => data <= "000000";
				when "001010101000000000" => data <= "000000";
				when "001010101000000001" => data <= "000000";
				when "001010101000000010" => data <= "000000";
				when "001010101000000011" => data <= "000000";
				when "001010101000000100" => data <= "000000";
				when "001010101000000101" => data <= "000000";
				when "001010101000000110" => data <= "000000";
				when "001010101000000111" => data <= "000000";
				when "001010101000001000" => data <= "000000";
				when "001010101000001001" => data <= "000000";
				when "001010101000001010" => data <= "000000";
				when "001010101000001011" => data <= "000000";
				when "001010101000001100" => data <= "000000";
				when "001010101000001101" => data <= "000000";
				when "001010101000001110" => data <= "000000";
				when "001010101000001111" => data <= "000000";
				when "001010101000010000" => data <= "000000";
				when "001010101000010001" => data <= "000000";
				when "001010101000010010" => data <= "000000";
				when "001010101000010011" => data <= "000000";
				when "001010101000010100" => data <= "000000";
				when "001010101000010101" => data <= "000000";
				when "001010101000010110" => data <= "000000";
				when "001010101000010111" => data <= "000000";
				when "001010101000011000" => data <= "000000";
				when "001010101000011001" => data <= "000000";
				when "001010101000011010" => data <= "000000";
				when "001010101000011011" => data <= "000000";
				when "001010101000011100" => data <= "000000";
				when "001010101000011101" => data <= "000000";
				when "001010101000011110" => data <= "000000";
				when "001010101000011111" => data <= "000000";
				when "001010101000100000" => data <= "000000";
				when "001010101000100001" => data <= "000000";
				when "001010101000100010" => data <= "000000";
				when "001010101000100011" => data <= "000000";
				when "001010101000100100" => data <= "000000";
				when "001010101000100101" => data <= "000000";
				when "001010101000100110" => data <= "000000";
				when "001010101000100111" => data <= "000000";
				when "001010101000101000" => data <= "000000";
				when "001010101000101001" => data <= "000000";
				when "001010101000101010" => data <= "000000";
				when "001010101000101011" => data <= "000000";
				when "001010101000101100" => data <= "000000";
				when "001010101000101101" => data <= "000000";
				when "001010101000101110" => data <= "000000";
				when "001010101000101111" => data <= "000000";
				when "001010101000110000" => data <= "000000";
				when "001010101000110001" => data <= "000000";
				when "001010101000110010" => data <= "000000";
				when "001010101000110011" => data <= "000000";
				when "001010101000110100" => data <= "000000";
				when "001010101000110101" => data <= "000000";
				when "001010101000110110" => data <= "000000";
				when "001010101000110111" => data <= "000000";
				when "001010101000111000" => data <= "000000";
				when "001010101000111001" => data <= "000000";
				when "001010101000111010" => data <= "000000";
				when "001010101000111011" => data <= "000000";
				when "001010101000111100" => data <= "000000";
				when "001010101000111101" => data <= "000000";
				when "001010101000111110" => data <= "000000";
				when "001010101000111111" => data <= "000000";
				when "001010101001000000" => data <= "000000";
				when "001010101001000001" => data <= "000000";
				when "001010101001000010" => data <= "000000";
				when "001010101001000011" => data <= "000000";
				when "001010101001000100" => data <= "000000";
				when "001010101001000101" => data <= "000000";
				when "001010101001000110" => data <= "000000";
				when "001010101001000111" => data <= "000000";
				when "001010101001001000" => data <= "000000";
				when "001010101001001001" => data <= "000000";
				when "001010101001001010" => data <= "000000";
				when "001010101001001011" => data <= "000000";
				when "001010101001001100" => data <= "000000";
				when "001010101001001101" => data <= "000000";
				when "001010101001001110" => data <= "000000";
				when "001010101001001111" => data <= "000000";
				when "001010101001010000" => data <= "000000";
				when "001010101001010001" => data <= "000000";
				when "001010101001010010" => data <= "000000";
				when "001010101001010011" => data <= "000000";
				when "001010101001010100" => data <= "000000";
				when "001010101001010101" => data <= "000000";
				when "001010101001010110" => data <= "000000";
				when "001010101001010111" => data <= "000000";
				when "001010101001011000" => data <= "000000";
				when "001010101001011001" => data <= "000000";
				when "001010101001011010" => data <= "000000";
				when "001010101001011011" => data <= "000000";
				when "001010101001011100" => data <= "000000";
				when "001010101001011101" => data <= "000000";
				when "001010101001011110" => data <= "000000";
				when "001010101001011111" => data <= "000000";
				when "001010101001100000" => data <= "000000";
				when "001010101001100001" => data <= "000000";
				when "001010101001100010" => data <= "000000";
				when "001010101001100011" => data <= "000000";
				when "001010101001100100" => data <= "000000";
				when "001010101001100101" => data <= "000000";
				when "001010101001100110" => data <= "000000";
				when "001010101001100111" => data <= "000000";
				when "001010101001101000" => data <= "000000";
				when "001010101001101001" => data <= "000000";
				when "001010101001101010" => data <= "000000";
				when "001010101001101011" => data <= "000000";
				when "001010101001101100" => data <= "000000";
				when "001010101001101101" => data <= "000000";
				when "001010101001101110" => data <= "000000";
				when "001010101001101111" => data <= "000000";
				when "001010101001110000" => data <= "000000";
				when "001010101001110001" => data <= "000000";
				when "001010101001110010" => data <= "000000";
				when "001010101001110011" => data <= "000000";
				when "001010101001110100" => data <= "000000";
				when "001010101001110101" => data <= "000000";
				when "001010101001110110" => data <= "000000";
				when "001010101001110111" => data <= "000000";
				when "001010101001111000" => data <= "000000";
				when "001010101001111001" => data <= "000000";
				when "001010101001111010" => data <= "000000";
				when "001010101001111011" => data <= "000000";
				when "001010101001111100" => data <= "000000";
				when "001010101001111101" => data <= "000000";
				when "001010101001111110" => data <= "000000";
				when "001010101001111111" => data <= "000000";
				when "001010101010000000" => data <= "000000";
				when "001010101010000001" => data <= "000000";
				when "001010101010000010" => data <= "000000";
				when "001010101010000011" => data <= "000000";
				when "001010101010000100" => data <= "000000";
				when "001010101010000101" => data <= "000000";
				when "001010101010000110" => data <= "000000";
				when "001010101010000111" => data <= "000000";
				when "001010101010001000" => data <= "000000";
				when "001010101010001001" => data <= "000000";
				when "001010101010001010" => data <= "000000";
				when "001010101010001011" => data <= "000000";
				when "001010101010001100" => data <= "000000";
				when "001010101010001101" => data <= "000000";
				when "001010101010001110" => data <= "000000";
				when "001010101010001111" => data <= "000000";
				when "001010101010010000" => data <= "000000";
				when "001010101010010001" => data <= "000000";
				when "001010101010010010" => data <= "000000";
				when "001010101010010011" => data <= "000000";
				when "001010101010010100" => data <= "000000";
				when "001010101010010101" => data <= "000000";
				when "001010101010010110" => data <= "000000";
				when "001010101010010111" => data <= "000000";
				when "001010101010011000" => data <= "000000";
				when "001010101010011001" => data <= "000000";
				when "001010101010011010" => data <= "000000";
				when "001010101010011011" => data <= "000000";
				when "001010101010011100" => data <= "000000";
				when "001010101010011101" => data <= "000000";
				when "001010101010011110" => data <= "000000";
				when "001010101010011111" => data <= "000000";
				when "001010110000000000" => data <= "000000";
				when "001010110000000001" => data <= "000000";
				when "001010110000000010" => data <= "000000";
				when "001010110000000011" => data <= "000000";
				when "001010110000000100" => data <= "000000";
				when "001010110000000101" => data <= "000000";
				when "001010110000000110" => data <= "000000";
				when "001010110000000111" => data <= "000000";
				when "001010110000001000" => data <= "000000";
				when "001010110000001001" => data <= "000000";
				when "001010110000001010" => data <= "000000";
				when "001010110000001011" => data <= "000000";
				when "001010110000001100" => data <= "000000";
				when "001010110000001101" => data <= "000000";
				when "001010110000001110" => data <= "000000";
				when "001010110000001111" => data <= "000000";
				when "001010110000010000" => data <= "000000";
				when "001010110000010001" => data <= "000000";
				when "001010110000010010" => data <= "000000";
				when "001010110000010011" => data <= "000000";
				when "001010110000010100" => data <= "000000";
				when "001010110000010101" => data <= "000000";
				when "001010110000010110" => data <= "000000";
				when "001010110000010111" => data <= "000000";
				when "001010110000011000" => data <= "000000";
				when "001010110000011001" => data <= "000000";
				when "001010110000011010" => data <= "000000";
				when "001010110000011011" => data <= "000000";
				when "001010110000011100" => data <= "000000";
				when "001010110000011101" => data <= "000000";
				when "001010110000011110" => data <= "000000";
				when "001010110000011111" => data <= "000000";
				when "001010110000100000" => data <= "000000";
				when "001010110000100001" => data <= "000000";
				when "001010110000100010" => data <= "000000";
				when "001010110000100011" => data <= "000000";
				when "001010110000100100" => data <= "000000";
				when "001010110000100101" => data <= "000000";
				when "001010110000100110" => data <= "000000";
				when "001010110000100111" => data <= "000000";
				when "001010110000101000" => data <= "000000";
				when "001010110000101001" => data <= "000000";
				when "001010110000101010" => data <= "000000";
				when "001010110000101011" => data <= "000000";
				when "001010110000101100" => data <= "000000";
				when "001010110000101101" => data <= "000000";
				when "001010110000101110" => data <= "000000";
				when "001010110000101111" => data <= "000000";
				when "001010110000110000" => data <= "000000";
				when "001010110000110001" => data <= "000000";
				when "001010110000110010" => data <= "000000";
				when "001010110000110011" => data <= "000000";
				when "001010110000110100" => data <= "000000";
				when "001010110000110101" => data <= "000000";
				when "001010110000110110" => data <= "000000";
				when "001010110000110111" => data <= "000000";
				when "001010110000111000" => data <= "000000";
				when "001010110000111001" => data <= "000000";
				when "001010110000111010" => data <= "000000";
				when "001010110000111011" => data <= "000000";
				when "001010110000111100" => data <= "000000";
				when "001010110000111101" => data <= "000000";
				when "001010110000111110" => data <= "000000";
				when "001010110000111111" => data <= "000000";
				when "001010110001000000" => data <= "000000";
				when "001010110001000001" => data <= "000000";
				when "001010110001000010" => data <= "000000";
				when "001010110001000011" => data <= "000000";
				when "001010110001000100" => data <= "000000";
				when "001010110001000101" => data <= "000000";
				when "001010110001000110" => data <= "000000";
				when "001010110001000111" => data <= "000000";
				when "001010110001001000" => data <= "000000";
				when "001010110001001001" => data <= "000000";
				when "001010110001001010" => data <= "000000";
				when "001010110001001011" => data <= "000000";
				when "001010110001001100" => data <= "000000";
				when "001010110001001101" => data <= "000000";
				when "001010110001001110" => data <= "000000";
				when "001010110001001111" => data <= "000000";
				when "001010110001010000" => data <= "000000";
				when "001010110001010001" => data <= "000000";
				when "001010110001010010" => data <= "000000";
				when "001010110001010011" => data <= "000000";
				when "001010110001010100" => data <= "000000";
				when "001010110001010101" => data <= "000000";
				when "001010110001010110" => data <= "000000";
				when "001010110001010111" => data <= "000000";
				when "001010110001011000" => data <= "000000";
				when "001010110001011001" => data <= "000000";
				when "001010110001011010" => data <= "000000";
				when "001010110001011011" => data <= "000000";
				when "001010110001011100" => data <= "000000";
				when "001010110001011101" => data <= "000000";
				when "001010110001011110" => data <= "000000";
				when "001010110001011111" => data <= "000000";
				when "001010110001100000" => data <= "000000";
				when "001010110001100001" => data <= "000000";
				when "001010110001100010" => data <= "000000";
				when "001010110001100011" => data <= "000000";
				when "001010110001100100" => data <= "000000";
				when "001010110001100101" => data <= "000000";
				when "001010110001100110" => data <= "000000";
				when "001010110001100111" => data <= "000000";
				when "001010110001101000" => data <= "000000";
				when "001010110001101001" => data <= "000000";
				when "001010110001101010" => data <= "000000";
				when "001010110001101011" => data <= "000000";
				when "001010110001101100" => data <= "000000";
				when "001010110001101101" => data <= "000000";
				when "001010110001101110" => data <= "000000";
				when "001010110001101111" => data <= "000000";
				when "001010110001110000" => data <= "000000";
				when "001010110001110001" => data <= "000000";
				when "001010110001110010" => data <= "000000";
				when "001010110001110011" => data <= "000000";
				when "001010110001110100" => data <= "000000";
				when "001010110001110101" => data <= "000000";
				when "001010110001110110" => data <= "000000";
				when "001010110001110111" => data <= "000000";
				when "001010110001111000" => data <= "000000";
				when "001010110001111001" => data <= "000000";
				when "001010110001111010" => data <= "000000";
				when "001010110001111011" => data <= "000000";
				when "001010110001111100" => data <= "000000";
				when "001010110001111101" => data <= "000000";
				when "001010110001111110" => data <= "000000";
				when "001010110001111111" => data <= "000000";
				when "001010110010000000" => data <= "000000";
				when "001010110010000001" => data <= "000000";
				when "001010110010000010" => data <= "000000";
				when "001010110010000011" => data <= "000000";
				when "001010110010000100" => data <= "000000";
				when "001010110010000101" => data <= "000000";
				when "001010110010000110" => data <= "000000";
				when "001010110010000111" => data <= "000000";
				when "001010110010001000" => data <= "000000";
				when "001010110010001001" => data <= "000000";
				when "001010110010001010" => data <= "000000";
				when "001010110010001011" => data <= "000000";
				when "001010110010001100" => data <= "000000";
				when "001010110010001101" => data <= "000000";
				when "001010110010001110" => data <= "000000";
				when "001010110010001111" => data <= "000000";
				when "001010110010010000" => data <= "000000";
				when "001010110010010001" => data <= "000000";
				when "001010110010010010" => data <= "000000";
				when "001010110010010011" => data <= "000000";
				when "001010110010010100" => data <= "000000";
				when "001010110010010101" => data <= "000000";
				when "001010110010010110" => data <= "000000";
				when "001010110010010111" => data <= "000000";
				when "001010110010011000" => data <= "000000";
				when "001010110010011001" => data <= "000000";
				when "001010110010011010" => data <= "000000";
				when "001010110010011011" => data <= "000000";
				when "001010110010011100" => data <= "000000";
				when "001010110010011101" => data <= "000000";
				when "001010110010011110" => data <= "000000";
				when "001010110010011111" => data <= "000000";
				when "001010111000000000" => data <= "000000";
				when "001010111000000001" => data <= "000000";
				when "001010111000000010" => data <= "000000";
				when "001010111000000011" => data <= "000000";
				when "001010111000000100" => data <= "000000";
				when "001010111000000101" => data <= "000000";
				when "001010111000000110" => data <= "000000";
				when "001010111000000111" => data <= "000000";
				when "001010111000001000" => data <= "000000";
				when "001010111000001001" => data <= "000000";
				when "001010111000001010" => data <= "000000";
				when "001010111000001011" => data <= "000000";
				when "001010111000001100" => data <= "000000";
				when "001010111000001101" => data <= "000000";
				when "001010111000001110" => data <= "000000";
				when "001010111000001111" => data <= "000000";
				when "001010111000010000" => data <= "000000";
				when "001010111000010001" => data <= "000000";
				when "001010111000010010" => data <= "000000";
				when "001010111000010011" => data <= "000000";
				when "001010111000010100" => data <= "000000";
				when "001010111000010101" => data <= "000000";
				when "001010111000010110" => data <= "000000";
				when "001010111000010111" => data <= "000000";
				when "001010111000011000" => data <= "000000";
				when "001010111000011001" => data <= "000000";
				when "001010111000011010" => data <= "000000";
				when "001010111000011011" => data <= "000000";
				when "001010111000011100" => data <= "000000";
				when "001010111000011101" => data <= "000000";
				when "001010111000011110" => data <= "000000";
				when "001010111000011111" => data <= "000000";
				when "001010111000100000" => data <= "000000";
				when "001010111000100001" => data <= "000000";
				when "001010111000100010" => data <= "000000";
				when "001010111000100011" => data <= "000000";
				when "001010111000100100" => data <= "000000";
				when "001010111000100101" => data <= "000000";
				when "001010111000100110" => data <= "000000";
				when "001010111000100111" => data <= "000000";
				when "001010111000101000" => data <= "000000";
				when "001010111000101001" => data <= "000000";
				when "001010111000101010" => data <= "000000";
				when "001010111000101011" => data <= "000000";
				when "001010111000101100" => data <= "000000";
				when "001010111000101101" => data <= "000000";
				when "001010111000101110" => data <= "000000";
				when "001010111000101111" => data <= "000000";
				when "001010111000110000" => data <= "000000";
				when "001010111000110001" => data <= "000000";
				when "001010111000110010" => data <= "000000";
				when "001010111000110011" => data <= "000000";
				when "001010111000110100" => data <= "000000";
				when "001010111000110101" => data <= "000000";
				when "001010111000110110" => data <= "000000";
				when "001010111000110111" => data <= "000000";
				when "001010111000111000" => data <= "000000";
				when "001010111000111001" => data <= "000000";
				when "001010111000111010" => data <= "000000";
				when "001010111000111011" => data <= "000000";
				when "001010111000111100" => data <= "000000";
				when "001010111000111101" => data <= "000000";
				when "001010111000111110" => data <= "000000";
				when "001010111000111111" => data <= "000000";
				when "001010111001000000" => data <= "000000";
				when "001010111001000001" => data <= "000000";
				when "001010111001000010" => data <= "000000";
				when "001010111001000011" => data <= "000000";
				when "001010111001000100" => data <= "000000";
				when "001010111001000101" => data <= "000000";
				when "001010111001000110" => data <= "000000";
				when "001010111001000111" => data <= "000000";
				when "001010111001001000" => data <= "000000";
				when "001010111001001001" => data <= "000000";
				when "001010111001001010" => data <= "000000";
				when "001010111001001011" => data <= "000000";
				when "001010111001001100" => data <= "000000";
				when "001010111001001101" => data <= "000000";
				when "001010111001001110" => data <= "000000";
				when "001010111001001111" => data <= "000000";
				when "001010111001010000" => data <= "000000";
				when "001010111001010001" => data <= "000000";
				when "001010111001010010" => data <= "000000";
				when "001010111001010011" => data <= "000000";
				when "001010111001010100" => data <= "000000";
				when "001010111001010101" => data <= "000000";
				when "001010111001010110" => data <= "000000";
				when "001010111001010111" => data <= "000000";
				when "001010111001011000" => data <= "000000";
				when "001010111001011001" => data <= "000000";
				when "001010111001011010" => data <= "000000";
				when "001010111001011011" => data <= "000000";
				when "001010111001011100" => data <= "000000";
				when "001010111001011101" => data <= "000000";
				when "001010111001011110" => data <= "000000";
				when "001010111001011111" => data <= "000000";
				when "001010111001100000" => data <= "000000";
				when "001010111001100001" => data <= "000000";
				when "001010111001100010" => data <= "000000";
				when "001010111001100011" => data <= "000000";
				when "001010111001100100" => data <= "000000";
				when "001010111001100101" => data <= "000000";
				when "001010111001100110" => data <= "000000";
				when "001010111001100111" => data <= "000000";
				when "001010111001101000" => data <= "000000";
				when "001010111001101001" => data <= "000000";
				when "001010111001101010" => data <= "000000";
				when "001010111001101011" => data <= "000000";
				when "001010111001101100" => data <= "000000";
				when "001010111001101101" => data <= "000000";
				when "001010111001101110" => data <= "000000";
				when "001010111001101111" => data <= "000000";
				when "001010111001110000" => data <= "000000";
				when "001010111001110001" => data <= "000000";
				when "001010111001110010" => data <= "000000";
				when "001010111001110011" => data <= "000000";
				when "001010111001110100" => data <= "000000";
				when "001010111001110101" => data <= "000000";
				when "001010111001110110" => data <= "000000";
				when "001010111001110111" => data <= "000000";
				when "001010111001111000" => data <= "000000";
				when "001010111001111001" => data <= "000000";
				when "001010111001111010" => data <= "000000";
				when "001010111001111011" => data <= "000000";
				when "001010111001111100" => data <= "000000";
				when "001010111001111101" => data <= "000000";
				when "001010111001111110" => data <= "000000";
				when "001010111001111111" => data <= "000000";
				when "001010111010000000" => data <= "000000";
				when "001010111010000001" => data <= "000000";
				when "001010111010000010" => data <= "000000";
				when "001010111010000011" => data <= "000000";
				when "001010111010000100" => data <= "000000";
				when "001010111010000101" => data <= "000000";
				when "001010111010000110" => data <= "000000";
				when "001010111010000111" => data <= "000000";
				when "001010111010001000" => data <= "000000";
				when "001010111010001001" => data <= "000000";
				when "001010111010001010" => data <= "000000";
				when "001010111010001011" => data <= "000000";
				when "001010111010001100" => data <= "000000";
				when "001010111010001101" => data <= "000000";
				when "001010111010001110" => data <= "000000";
				when "001010111010001111" => data <= "000000";
				when "001010111010010000" => data <= "000000";
				when "001010111010010001" => data <= "000000";
				when "001010111010010010" => data <= "000000";
				when "001010111010010011" => data <= "000000";
				when "001010111010010100" => data <= "000000";
				when "001010111010010101" => data <= "000000";
				when "001010111010010110" => data <= "000000";
				when "001010111010010111" => data <= "000000";
				when "001010111010011000" => data <= "000000";
				when "001010111010011001" => data <= "000000";
				when "001010111010011010" => data <= "000000";
				when "001010111010011011" => data <= "000000";
				when "001010111010011100" => data <= "000000";
				when "001010111010011101" => data <= "000000";
				when "001010111010011110" => data <= "000000";
				when "001010111010011111" => data <= "000000";
				when "001011000000000000" => data <= "000000";
				when "001011000000000001" => data <= "000000";
				when "001011000000000010" => data <= "000000";
				when "001011000000000011" => data <= "000000";
				when "001011000000000100" => data <= "000000";
				when "001011000000000101" => data <= "000000";
				when "001011000000000110" => data <= "000000";
				when "001011000000000111" => data <= "000000";
				when "001011000000001000" => data <= "000000";
				when "001011000000001001" => data <= "000000";
				when "001011000000001010" => data <= "000000";
				when "001011000000001011" => data <= "000000";
				when "001011000000001100" => data <= "000000";
				when "001011000000001101" => data <= "000000";
				when "001011000000001110" => data <= "000000";
				when "001011000000001111" => data <= "000000";
				when "001011000000010000" => data <= "000000";
				when "001011000000010001" => data <= "000000";
				when "001011000000010010" => data <= "000000";
				when "001011000000010011" => data <= "000000";
				when "001011000000010100" => data <= "000000";
				when "001011000000010101" => data <= "000000";
				when "001011000000010110" => data <= "000000";
				when "001011000000010111" => data <= "000000";
				when "001011000000011000" => data <= "000000";
				when "001011000000011001" => data <= "000000";
				when "001011000000011010" => data <= "000000";
				when "001011000000011011" => data <= "000000";
				when "001011000000011100" => data <= "000000";
				when "001011000000011101" => data <= "000000";
				when "001011000000011110" => data <= "000000";
				when "001011000000011111" => data <= "000000";
				when "001011000000100000" => data <= "000000";
				when "001011000000100001" => data <= "000000";
				when "001011000000100010" => data <= "000000";
				when "001011000000100011" => data <= "000000";
				when "001011000000100100" => data <= "000000";
				when "001011000000100101" => data <= "000000";
				when "001011000000100110" => data <= "000000";
				when "001011000000100111" => data <= "000000";
				when "001011000000101000" => data <= "000000";
				when "001011000000101001" => data <= "000000";
				when "001011000000101010" => data <= "000000";
				when "001011000000101011" => data <= "000000";
				when "001011000000101100" => data <= "000000";
				when "001011000000101101" => data <= "000000";
				when "001011000000101110" => data <= "000000";
				when "001011000000101111" => data <= "000000";
				when "001011000000110000" => data <= "000000";
				when "001011000000110001" => data <= "000000";
				when "001011000000110010" => data <= "000000";
				when "001011000000110011" => data <= "000000";
				when "001011000000110100" => data <= "000000";
				when "001011000000110101" => data <= "000000";
				when "001011000000110110" => data <= "000000";
				when "001011000000110111" => data <= "000000";
				when "001011000000111000" => data <= "000000";
				when "001011000000111001" => data <= "000000";
				when "001011000000111010" => data <= "000000";
				when "001011000000111011" => data <= "000000";
				when "001011000000111100" => data <= "000000";
				when "001011000000111101" => data <= "000000";
				when "001011000000111110" => data <= "000000";
				when "001011000000111111" => data <= "000000";
				when "001011000001000000" => data <= "000000";
				when "001011000001000001" => data <= "000000";
				when "001011000001000010" => data <= "000000";
				when "001011000001000011" => data <= "000000";
				when "001011000001000100" => data <= "000000";
				when "001011000001000101" => data <= "000000";
				when "001011000001000110" => data <= "000000";
				when "001011000001000111" => data <= "000000";
				when "001011000001001000" => data <= "000000";
				when "001011000001001001" => data <= "000000";
				when "001011000001001010" => data <= "000000";
				when "001011000001001011" => data <= "000000";
				when "001011000001001100" => data <= "000000";
				when "001011000001001101" => data <= "000000";
				when "001011000001001110" => data <= "000000";
				when "001011000001001111" => data <= "000000";
				when "001011000001010000" => data <= "000000";
				when "001011000001010001" => data <= "000000";
				when "001011000001010010" => data <= "000000";
				when "001011000001010011" => data <= "000000";
				when "001011000001010100" => data <= "000000";
				when "001011000001010101" => data <= "000000";
				when "001011000001010110" => data <= "000000";
				when "001011000001010111" => data <= "000000";
				when "001011000001011000" => data <= "000000";
				when "001011000001011001" => data <= "000000";
				when "001011000001011010" => data <= "000000";
				when "001011000001011011" => data <= "000000";
				when "001011000001011100" => data <= "000000";
				when "001011000001011101" => data <= "000000";
				when "001011000001011110" => data <= "000000";
				when "001011000001011111" => data <= "000000";
				when "001011000001100000" => data <= "000000";
				when "001011000001100001" => data <= "000000";
				when "001011000001100010" => data <= "000000";
				when "001011000001100011" => data <= "000000";
				when "001011000001100100" => data <= "000000";
				when "001011000001100101" => data <= "000000";
				when "001011000001100110" => data <= "000000";
				when "001011000001100111" => data <= "000000";
				when "001011000001101000" => data <= "000000";
				when "001011000001101001" => data <= "000000";
				when "001011000001101010" => data <= "000000";
				when "001011000001101011" => data <= "000000";
				when "001011000001101100" => data <= "000000";
				when "001011000001101101" => data <= "000000";
				when "001011000001101110" => data <= "000000";
				when "001011000001101111" => data <= "000000";
				when "001011000001110000" => data <= "000000";
				when "001011000001110001" => data <= "000000";
				when "001011000001110010" => data <= "000000";
				when "001011000001110011" => data <= "000000";
				when "001011000001110100" => data <= "000000";
				when "001011000001110101" => data <= "000000";
				when "001011000001110110" => data <= "000000";
				when "001011000001110111" => data <= "000000";
				when "001011000001111000" => data <= "000000";
				when "001011000001111001" => data <= "000000";
				when "001011000001111010" => data <= "000000";
				when "001011000001111011" => data <= "000000";
				when "001011000001111100" => data <= "000000";
				when "001011000001111101" => data <= "000000";
				when "001011000001111110" => data <= "000000";
				when "001011000001111111" => data <= "000000";
				when "001011000010000000" => data <= "000000";
				when "001011000010000001" => data <= "000000";
				when "001011000010000010" => data <= "000000";
				when "001011000010000011" => data <= "000000";
				when "001011000010000100" => data <= "000000";
				when "001011000010000101" => data <= "000000";
				when "001011000010000110" => data <= "000000";
				when "001011000010000111" => data <= "000000";
				when "001011000010001000" => data <= "000000";
				when "001011000010001001" => data <= "000000";
				when "001011000010001010" => data <= "000000";
				when "001011000010001011" => data <= "000000";
				when "001011000010001100" => data <= "000000";
				when "001011000010001101" => data <= "000000";
				when "001011000010001110" => data <= "000000";
				when "001011000010001111" => data <= "000000";
				when "001011000010010000" => data <= "000000";
				when "001011000010010001" => data <= "000000";
				when "001011000010010010" => data <= "000000";
				when "001011000010010011" => data <= "000000";
				when "001011000010010100" => data <= "000000";
				when "001011000010010101" => data <= "000000";
				when "001011000010010110" => data <= "000000";
				when "001011000010010111" => data <= "000000";
				when "001011000010011000" => data <= "000000";
				when "001011000010011001" => data <= "000000";
				when "001011000010011010" => data <= "000000";
				when "001011000010011011" => data <= "000000";
				when "001011000010011100" => data <= "000000";
				when "001011000010011101" => data <= "000000";
				when "001011000010011110" => data <= "000000";
				when "001011000010011111" => data <= "000000";
				when "001011001000000000" => data <= "000000";
				when "001011001000000001" => data <= "000000";
				when "001011001000000010" => data <= "000000";
				when "001011001000000011" => data <= "000000";
				when "001011001000000100" => data <= "000000";
				when "001011001000000101" => data <= "000000";
				when "001011001000000110" => data <= "000000";
				when "001011001000000111" => data <= "000000";
				when "001011001000001000" => data <= "000000";
				when "001011001000001001" => data <= "000000";
				when "001011001000001010" => data <= "000000";
				when "001011001000001011" => data <= "000000";
				when "001011001000001100" => data <= "000000";
				when "001011001000001101" => data <= "000000";
				when "001011001000001110" => data <= "000000";
				when "001011001000001111" => data <= "000000";
				when "001011001000010000" => data <= "000000";
				when "001011001000010001" => data <= "000000";
				when "001011001000010010" => data <= "000000";
				when "001011001000010011" => data <= "000000";
				when "001011001000010100" => data <= "000000";
				when "001011001000010101" => data <= "000000";
				when "001011001000010110" => data <= "000000";
				when "001011001000010111" => data <= "000000";
				when "001011001000011000" => data <= "000000";
				when "001011001000011001" => data <= "000000";
				when "001011001000011010" => data <= "000000";
				when "001011001000011011" => data <= "000000";
				when "001011001000011100" => data <= "000000";
				when "001011001000011101" => data <= "000000";
				when "001011001000011110" => data <= "000000";
				when "001011001000011111" => data <= "000000";
				when "001011001000100000" => data <= "000000";
				when "001011001000100001" => data <= "000000";
				when "001011001000100010" => data <= "000000";
				when "001011001000100011" => data <= "000000";
				when "001011001000100100" => data <= "000000";
				when "001011001000100101" => data <= "000000";
				when "001011001000100110" => data <= "000000";
				when "001011001000100111" => data <= "000000";
				when "001011001000101000" => data <= "000000";
				when "001011001000101001" => data <= "000000";
				when "001011001000101010" => data <= "000000";
				when "001011001000101011" => data <= "000000";
				when "001011001000101100" => data <= "000000";
				when "001011001000101101" => data <= "000000";
				when "001011001000101110" => data <= "000000";
				when "001011001000101111" => data <= "000000";
				when "001011001000110000" => data <= "000000";
				when "001011001000110001" => data <= "000000";
				when "001011001000110010" => data <= "000000";
				when "001011001000110011" => data <= "000000";
				when "001011001000110100" => data <= "000000";
				when "001011001000110101" => data <= "000000";
				when "001011001000110110" => data <= "000000";
				when "001011001000110111" => data <= "000000";
				when "001011001000111000" => data <= "000000";
				when "001011001000111001" => data <= "000000";
				when "001011001000111010" => data <= "000000";
				when "001011001000111011" => data <= "000000";
				when "001011001000111100" => data <= "000000";
				when "001011001000111101" => data <= "000000";
				when "001011001000111110" => data <= "000000";
				when "001011001000111111" => data <= "000000";
				when "001011001001000000" => data <= "000000";
				when "001011001001000001" => data <= "000000";
				when "001011001001000010" => data <= "000000";
				when "001011001001000011" => data <= "000000";
				when "001011001001000100" => data <= "000000";
				when "001011001001000101" => data <= "000000";
				when "001011001001000110" => data <= "000000";
				when "001011001001000111" => data <= "000000";
				when "001011001001001000" => data <= "000000";
				when "001011001001001001" => data <= "000000";
				when "001011001001001010" => data <= "000000";
				when "001011001001001011" => data <= "000000";
				when "001011001001001100" => data <= "000000";
				when "001011001001001101" => data <= "000000";
				when "001011001001001110" => data <= "000000";
				when "001011001001001111" => data <= "000000";
				when "001011001001010000" => data <= "000000";
				when "001011001001010001" => data <= "000000";
				when "001011001001010010" => data <= "000000";
				when "001011001001010011" => data <= "000000";
				when "001011001001010100" => data <= "000000";
				when "001011001001010101" => data <= "000000";
				when "001011001001010110" => data <= "000000";
				when "001011001001010111" => data <= "000000";
				when "001011001001011000" => data <= "000000";
				when "001011001001011001" => data <= "000000";
				when "001011001001011010" => data <= "000000";
				when "001011001001011011" => data <= "000000";
				when "001011001001011100" => data <= "000000";
				when "001011001001011101" => data <= "000000";
				when "001011001001011110" => data <= "000000";
				when "001011001001011111" => data <= "000000";
				when "001011001001100000" => data <= "000000";
				when "001011001001100001" => data <= "000000";
				when "001011001001100010" => data <= "000000";
				when "001011001001100011" => data <= "000000";
				when "001011001001100100" => data <= "000000";
				when "001011001001100101" => data <= "000000";
				when "001011001001100110" => data <= "000000";
				when "001011001001100111" => data <= "000000";
				when "001011001001101000" => data <= "000000";
				when "001011001001101001" => data <= "000000";
				when "001011001001101010" => data <= "000000";
				when "001011001001101011" => data <= "000000";
				when "001011001001101100" => data <= "000000";
				when "001011001001101101" => data <= "000000";
				when "001011001001101110" => data <= "000000";
				when "001011001001101111" => data <= "000000";
				when "001011001001110000" => data <= "000000";
				when "001011001001110001" => data <= "000000";
				when "001011001001110010" => data <= "000000";
				when "001011001001110011" => data <= "000000";
				when "001011001001110100" => data <= "000000";
				when "001011001001110101" => data <= "000000";
				when "001011001001110110" => data <= "000000";
				when "001011001001110111" => data <= "000000";
				when "001011001001111000" => data <= "000000";
				when "001011001001111001" => data <= "000000";
				when "001011001001111010" => data <= "000000";
				when "001011001001111011" => data <= "000000";
				when "001011001001111100" => data <= "000000";
				when "001011001001111101" => data <= "000000";
				when "001011001001111110" => data <= "000000";
				when "001011001001111111" => data <= "000000";
				when "001011001010000000" => data <= "000000";
				when "001011001010000001" => data <= "000000";
				when "001011001010000010" => data <= "000000";
				when "001011001010000011" => data <= "000000";
				when "001011001010000100" => data <= "000000";
				when "001011001010000101" => data <= "000000";
				when "001011001010000110" => data <= "000000";
				when "001011001010000111" => data <= "000000";
				when "001011001010001000" => data <= "000000";
				when "001011001010001001" => data <= "000000";
				when "001011001010001010" => data <= "000000";
				when "001011001010001011" => data <= "000000";
				when "001011001010001100" => data <= "000000";
				when "001011001010001101" => data <= "000000";
				when "001011001010001110" => data <= "000000";
				when "001011001010001111" => data <= "000000";
				when "001011001010010000" => data <= "000000";
				when "001011001010010001" => data <= "000000";
				when "001011001010010010" => data <= "000000";
				when "001011001010010011" => data <= "000000";
				when "001011001010010100" => data <= "000000";
				when "001011001010010101" => data <= "000000";
				when "001011001010010110" => data <= "000000";
				when "001011001010010111" => data <= "000000";
				when "001011001010011000" => data <= "000000";
				when "001011001010011001" => data <= "000000";
				when "001011001010011010" => data <= "000000";
				when "001011001010011011" => data <= "000000";
				when "001011001010011100" => data <= "000000";
				when "001011001010011101" => data <= "000000";
				when "001011001010011110" => data <= "000000";
				when "001011001010011111" => data <= "000000";
				when "001011010000000000" => data <= "000000";
				when "001011010000000001" => data <= "000000";
				when "001011010000000010" => data <= "000000";
				when "001011010000000011" => data <= "000000";
				when "001011010000000100" => data <= "000000";
				when "001011010000000101" => data <= "000000";
				when "001011010000000110" => data <= "000000";
				when "001011010000000111" => data <= "000000";
				when "001011010000001000" => data <= "000000";
				when "001011010000001001" => data <= "000000";
				when "001011010000001010" => data <= "000000";
				when "001011010000001011" => data <= "000000";
				when "001011010000001100" => data <= "000000";
				when "001011010000001101" => data <= "000000";
				when "001011010000001110" => data <= "000000";
				when "001011010000001111" => data <= "000000";
				when "001011010000010000" => data <= "000000";
				when "001011010000010001" => data <= "000000";
				when "001011010000010010" => data <= "000000";
				when "001011010000010011" => data <= "000000";
				when "001011010000010100" => data <= "000000";
				when "001011010000010101" => data <= "000000";
				when "001011010000010110" => data <= "000000";
				when "001011010000010111" => data <= "000000";
				when "001011010000011000" => data <= "000000";
				when "001011010000011001" => data <= "000000";
				when "001011010000011010" => data <= "000000";
				when "001011010000011011" => data <= "000000";
				when "001011010000011100" => data <= "000000";
				when "001011010000011101" => data <= "000000";
				when "001011010000011110" => data <= "000000";
				when "001011010000011111" => data <= "000000";
				when "001011010000100000" => data <= "000000";
				when "001011010000100001" => data <= "000000";
				when "001011010000100010" => data <= "000000";
				when "001011010000100011" => data <= "000000";
				when "001011010000100100" => data <= "000000";
				when "001011010000100101" => data <= "000000";
				when "001011010000100110" => data <= "000000";
				when "001011010000100111" => data <= "000000";
				when "001011010000101000" => data <= "000000";
				when "001011010000101001" => data <= "000000";
				when "001011010000101010" => data <= "000000";
				when "001011010000101011" => data <= "000000";
				when "001011010000101100" => data <= "000000";
				when "001011010000101101" => data <= "000000";
				when "001011010000101110" => data <= "000000";
				when "001011010000101111" => data <= "000000";
				when "001011010000110000" => data <= "000000";
				when "001011010000110001" => data <= "000000";
				when "001011010000110010" => data <= "000000";
				when "001011010000110011" => data <= "000000";
				when "001011010000110100" => data <= "000000";
				when "001011010000110101" => data <= "000000";
				when "001011010000110110" => data <= "000000";
				when "001011010000110111" => data <= "000000";
				when "001011010000111000" => data <= "000000";
				when "001011010000111001" => data <= "000000";
				when "001011010000111010" => data <= "000000";
				when "001011010000111011" => data <= "000000";
				when "001011010000111100" => data <= "000000";
				when "001011010000111101" => data <= "000000";
				when "001011010000111110" => data <= "000000";
				when "001011010000111111" => data <= "000000";
				when "001011010001000000" => data <= "000000";
				when "001011010001000001" => data <= "000000";
				when "001011010001000010" => data <= "000000";
				when "001011010001000011" => data <= "000000";
				when "001011010001000100" => data <= "000000";
				when "001011010001000101" => data <= "000000";
				when "001011010001000110" => data <= "000000";
				when "001011010001000111" => data <= "000000";
				when "001011010001001000" => data <= "000000";
				when "001011010001001001" => data <= "000000";
				when "001011010001001010" => data <= "000000";
				when "001011010001001011" => data <= "000000";
				when "001011010001001100" => data <= "000000";
				when "001011010001001101" => data <= "000000";
				when "001011010001001110" => data <= "000000";
				when "001011010001001111" => data <= "000000";
				when "001011010001010000" => data <= "000000";
				when "001011010001010001" => data <= "000000";
				when "001011010001010010" => data <= "000000";
				when "001011010001010011" => data <= "000000";
				when "001011010001010100" => data <= "000000";
				when "001011010001010101" => data <= "000000";
				when "001011010001010110" => data <= "000000";
				when "001011010001010111" => data <= "000000";
				when "001011010001011000" => data <= "000000";
				when "001011010001011001" => data <= "000000";
				when "001011010001011010" => data <= "000000";
				when "001011010001011011" => data <= "000000";
				when "001011010001011100" => data <= "000000";
				when "001011010001011101" => data <= "000000";
				when "001011010001011110" => data <= "000000";
				when "001011010001011111" => data <= "000000";
				when "001011010001100000" => data <= "000000";
				when "001011010001100001" => data <= "000000";
				when "001011010001100010" => data <= "000000";
				when "001011010001100011" => data <= "000000";
				when "001011010001100100" => data <= "000000";
				when "001011010001100101" => data <= "000000";
				when "001011010001100110" => data <= "000000";
				when "001011010001100111" => data <= "000000";
				when "001011010001101000" => data <= "000000";
				when "001011010001101001" => data <= "000000";
				when "001011010001101010" => data <= "000000";
				when "001011010001101011" => data <= "000000";
				when "001011010001101100" => data <= "000000";
				when "001011010001101101" => data <= "000000";
				when "001011010001101110" => data <= "000000";
				when "001011010001101111" => data <= "000000";
				when "001011010001110000" => data <= "000000";
				when "001011010001110001" => data <= "000000";
				when "001011010001110010" => data <= "000000";
				when "001011010001110011" => data <= "000000";
				when "001011010001110100" => data <= "000000";
				when "001011010001110101" => data <= "000000";
				when "001011010001110110" => data <= "000000";
				when "001011010001110111" => data <= "000000";
				when "001011010001111000" => data <= "000000";
				when "001011010001111001" => data <= "000000";
				when "001011010001111010" => data <= "000000";
				when "001011010001111011" => data <= "000000";
				when "001011010001111100" => data <= "000000";
				when "001011010001111101" => data <= "000000";
				when "001011010001111110" => data <= "000000";
				when "001011010001111111" => data <= "000000";
				when "001011010010000000" => data <= "000000";
				when "001011010010000001" => data <= "000000";
				when "001011010010000010" => data <= "000000";
				when "001011010010000011" => data <= "000000";
				when "001011010010000100" => data <= "000000";
				when "001011010010000101" => data <= "000000";
				when "001011010010000110" => data <= "000000";
				when "001011010010000111" => data <= "000000";
				when "001011010010001000" => data <= "000000";
				when "001011010010001001" => data <= "000000";
				when "001011010010001010" => data <= "000000";
				when "001011010010001011" => data <= "000000";
				when "001011010010001100" => data <= "000000";
				when "001011010010001101" => data <= "000000";
				when "001011010010001110" => data <= "000000";
				when "001011010010001111" => data <= "000000";
				when "001011010010010000" => data <= "000000";
				when "001011010010010001" => data <= "000000";
				when "001011010010010010" => data <= "000000";
				when "001011010010010011" => data <= "000000";
				when "001011010010010100" => data <= "000000";
				when "001011010010010101" => data <= "000000";
				when "001011010010010110" => data <= "000000";
				when "001011010010010111" => data <= "000000";
				when "001011010010011000" => data <= "000000";
				when "001011010010011001" => data <= "000000";
				when "001011010010011010" => data <= "000000";
				when "001011010010011011" => data <= "000000";
				when "001011010010011100" => data <= "000000";
				when "001011010010011101" => data <= "000000";
				when "001011010010011110" => data <= "000000";
				when "001011010010011111" => data <= "000000";
				when "001011011000000000" => data <= "000000";
				when "001011011000000001" => data <= "000000";
				when "001011011000000010" => data <= "000000";
				when "001011011000000011" => data <= "000000";
				when "001011011000000100" => data <= "000000";
				when "001011011000000101" => data <= "000000";
				when "001011011000000110" => data <= "000000";
				when "001011011000000111" => data <= "000000";
				when "001011011000001000" => data <= "000000";
				when "001011011000001001" => data <= "000000";
				when "001011011000001010" => data <= "000000";
				when "001011011000001011" => data <= "000000";
				when "001011011000001100" => data <= "000000";
				when "001011011000001101" => data <= "000000";
				when "001011011000001110" => data <= "000000";
				when "001011011000001111" => data <= "000000";
				when "001011011000010000" => data <= "000000";
				when "001011011000010001" => data <= "000000";
				when "001011011000010010" => data <= "000000";
				when "001011011000010011" => data <= "000000";
				when "001011011000010100" => data <= "000000";
				when "001011011000010101" => data <= "000000";
				when "001011011000010110" => data <= "000000";
				when "001011011000010111" => data <= "000000";
				when "001011011000011000" => data <= "000000";
				when "001011011000011001" => data <= "000000";
				when "001011011000011010" => data <= "000000";
				when "001011011000011011" => data <= "000000";
				when "001011011000011100" => data <= "000000";
				when "001011011000011101" => data <= "000000";
				when "001011011000011110" => data <= "000000";
				when "001011011000011111" => data <= "000000";
				when "001011011000100000" => data <= "000000";
				when "001011011000100001" => data <= "000000";
				when "001011011000100010" => data <= "000000";
				when "001011011000100011" => data <= "000000";
				when "001011011000100100" => data <= "000000";
				when "001011011000100101" => data <= "000000";
				when "001011011000100110" => data <= "000000";
				when "001011011000100111" => data <= "000000";
				when "001011011000101000" => data <= "000000";
				when "001011011000101001" => data <= "000000";
				when "001011011000101010" => data <= "000000";
				when "001011011000101011" => data <= "000000";
				when "001011011000101100" => data <= "000000";
				when "001011011000101101" => data <= "000000";
				when "001011011000101110" => data <= "000000";
				when "001011011000101111" => data <= "000000";
				when "001011011000110000" => data <= "000000";
				when "001011011000110001" => data <= "000000";
				when "001011011000110010" => data <= "000000";
				when "001011011000110011" => data <= "000000";
				when "001011011000110100" => data <= "000000";
				when "001011011000110101" => data <= "000000";
				when "001011011000110110" => data <= "000000";
				when "001011011000110111" => data <= "000000";
				when "001011011000111000" => data <= "000000";
				when "001011011000111001" => data <= "000000";
				when "001011011000111010" => data <= "000000";
				when "001011011000111011" => data <= "000000";
				when "001011011000111100" => data <= "000000";
				when "001011011000111101" => data <= "000000";
				when "001011011000111110" => data <= "000000";
				when "001011011000111111" => data <= "000000";
				when "001011011001000000" => data <= "000000";
				when "001011011001000001" => data <= "000000";
				when "001011011001000010" => data <= "000000";
				when "001011011001000011" => data <= "000000";
				when "001011011001000100" => data <= "000000";
				when "001011011001000101" => data <= "000000";
				when "001011011001000110" => data <= "000000";
				when "001011011001000111" => data <= "000000";
				when "001011011001001000" => data <= "000000";
				when "001011011001001001" => data <= "000000";
				when "001011011001001010" => data <= "000000";
				when "001011011001001011" => data <= "000000";
				when "001011011001001100" => data <= "000000";
				when "001011011001001101" => data <= "000000";
				when "001011011001001110" => data <= "000000";
				when "001011011001001111" => data <= "000000";
				when "001011011001010000" => data <= "000000";
				when "001011011001010001" => data <= "000000";
				when "001011011001010010" => data <= "000000";
				when "001011011001010011" => data <= "000000";
				when "001011011001010100" => data <= "000000";
				when "001011011001010101" => data <= "000000";
				when "001011011001010110" => data <= "000000";
				when "001011011001010111" => data <= "000000";
				when "001011011001011000" => data <= "000000";
				when "001011011001011001" => data <= "000000";
				when "001011011001011010" => data <= "000000";
				when "001011011001011011" => data <= "000000";
				when "001011011001011100" => data <= "000000";
				when "001011011001011101" => data <= "000000";
				when "001011011001011110" => data <= "000000";
				when "001011011001011111" => data <= "000000";
				when "001011011001100000" => data <= "000000";
				when "001011011001100001" => data <= "000000";
				when "001011011001100010" => data <= "000000";
				when "001011011001100011" => data <= "000000";
				when "001011011001100100" => data <= "000000";
				when "001011011001100101" => data <= "000000";
				when "001011011001100110" => data <= "000000";
				when "001011011001100111" => data <= "000000";
				when "001011011001101000" => data <= "000000";
				when "001011011001101001" => data <= "000000";
				when "001011011001101010" => data <= "000000";
				when "001011011001101011" => data <= "000000";
				when "001011011001101100" => data <= "000000";
				when "001011011001101101" => data <= "000000";
				when "001011011001101110" => data <= "000000";
				when "001011011001101111" => data <= "000000";
				when "001011011001110000" => data <= "000000";
				when "001011011001110001" => data <= "000000";
				when "001011011001110010" => data <= "000000";
				when "001011011001110011" => data <= "000000";
				when "001011011001110100" => data <= "000000";
				when "001011011001110101" => data <= "000000";
				when "001011011001110110" => data <= "000000";
				when "001011011001110111" => data <= "000000";
				when "001011011001111000" => data <= "000000";
				when "001011011001111001" => data <= "000000";
				when "001011011001111010" => data <= "000000";
				when "001011011001111011" => data <= "000000";
				when "001011011001111100" => data <= "000000";
				when "001011011001111101" => data <= "000000";
				when "001011011001111110" => data <= "000000";
				when "001011011001111111" => data <= "000000";
				when "001011011010000000" => data <= "000000";
				when "001011011010000001" => data <= "000000";
				when "001011011010000010" => data <= "000000";
				when "001011011010000011" => data <= "000000";
				when "001011011010000100" => data <= "000000";
				when "001011011010000101" => data <= "000000";
				when "001011011010000110" => data <= "000000";
				when "001011011010000111" => data <= "000000";
				when "001011011010001000" => data <= "000000";
				when "001011011010001001" => data <= "000000";
				when "001011011010001010" => data <= "000000";
				when "001011011010001011" => data <= "000000";
				when "001011011010001100" => data <= "000000";
				when "001011011010001101" => data <= "000000";
				when "001011011010001110" => data <= "000000";
				when "001011011010001111" => data <= "000000";
				when "001011011010010000" => data <= "000000";
				when "001011011010010001" => data <= "000000";
				when "001011011010010010" => data <= "000000";
				when "001011011010010011" => data <= "000000";
				when "001011011010010100" => data <= "000000";
				when "001011011010010101" => data <= "000000";
				when "001011011010010110" => data <= "000000";
				when "001011011010010111" => data <= "000000";
				when "001011011010011000" => data <= "000000";
				when "001011011010011001" => data <= "000000";
				when "001011011010011010" => data <= "000000";
				when "001011011010011011" => data <= "000000";
				when "001011011010011100" => data <= "000000";
				when "001011011010011101" => data <= "000000";
				when "001011011010011110" => data <= "000000";
				when "001011011010011111" => data <= "000000";
				when "001011100000000000" => data <= "000000";
				when "001011100000000001" => data <= "000000";
				when "001011100000000010" => data <= "000000";
				when "001011100000000011" => data <= "000000";
				when "001011100000000100" => data <= "000000";
				when "001011100000000101" => data <= "000000";
				when "001011100000000110" => data <= "000000";
				when "001011100000000111" => data <= "000000";
				when "001011100000001000" => data <= "000000";
				when "001011100000001001" => data <= "000000";
				when "001011100000001010" => data <= "000000";
				when "001011100000001011" => data <= "000000";
				when "001011100000001100" => data <= "000000";
				when "001011100000001101" => data <= "000000";
				when "001011100000001110" => data <= "000000";
				when "001011100000001111" => data <= "000000";
				when "001011100000010000" => data <= "000000";
				when "001011100000010001" => data <= "000000";
				when "001011100000010010" => data <= "000000";
				when "001011100000010011" => data <= "000000";
				when "001011100000010100" => data <= "000000";
				when "001011100000010101" => data <= "000000";
				when "001011100000010110" => data <= "000000";
				when "001011100000010111" => data <= "000000";
				when "001011100000011000" => data <= "000000";
				when "001011100000011001" => data <= "000000";
				when "001011100000011010" => data <= "000000";
				when "001011100000011011" => data <= "000000";
				when "001011100000011100" => data <= "000000";
				when "001011100000011101" => data <= "000000";
				when "001011100000011110" => data <= "000000";
				when "001011100000011111" => data <= "000000";
				when "001011100000100000" => data <= "000000";
				when "001011100000100001" => data <= "000000";
				when "001011100000100010" => data <= "000000";
				when "001011100000100011" => data <= "000000";
				when "001011100000100100" => data <= "000000";
				when "001011100000100101" => data <= "000000";
				when "001011100000100110" => data <= "000000";
				when "001011100000100111" => data <= "000000";
				when "001011100000101000" => data <= "000000";
				when "001011100000101001" => data <= "000000";
				when "001011100000101010" => data <= "000000";
				when "001011100000101011" => data <= "000000";
				when "001011100000101100" => data <= "000000";
				when "001011100000101101" => data <= "000000";
				when "001011100000101110" => data <= "000000";
				when "001011100000101111" => data <= "000000";
				when "001011100000110000" => data <= "000000";
				when "001011100000110001" => data <= "000000";
				when "001011100000110010" => data <= "000000";
				when "001011100000110011" => data <= "000000";
				when "001011100000110100" => data <= "000000";
				when "001011100000110101" => data <= "000000";
				when "001011100000110110" => data <= "000000";
				when "001011100000110111" => data <= "000000";
				when "001011100000111000" => data <= "000000";
				when "001011100000111001" => data <= "000000";
				when "001011100000111010" => data <= "000000";
				when "001011100000111011" => data <= "000000";
				when "001011100000111100" => data <= "000000";
				when "001011100000111101" => data <= "000000";
				when "001011100000111110" => data <= "000000";
				when "001011100000111111" => data <= "000000";
				when "001011100001000000" => data <= "000000";
				when "001011100001000001" => data <= "000000";
				when "001011100001000010" => data <= "000000";
				when "001011100001000011" => data <= "000000";
				when "001011100001000100" => data <= "000000";
				when "001011100001000101" => data <= "000000";
				when "001011100001000110" => data <= "000000";
				when "001011100001000111" => data <= "000000";
				when "001011100001001000" => data <= "000000";
				when "001011100001001001" => data <= "000000";
				when "001011100001001010" => data <= "000000";
				when "001011100001001011" => data <= "000000";
				when "001011100001001100" => data <= "000000";
				when "001011100001001101" => data <= "000000";
				when "001011100001001110" => data <= "000000";
				when "001011100001001111" => data <= "000000";
				when "001011100001010000" => data <= "000000";
				when "001011100001010001" => data <= "000000";
				when "001011100001010010" => data <= "000000";
				when "001011100001010011" => data <= "000000";
				when "001011100001010100" => data <= "000000";
				when "001011100001010101" => data <= "000000";
				when "001011100001010110" => data <= "000000";
				when "001011100001010111" => data <= "000000";
				when "001011100001011000" => data <= "000000";
				when "001011100001011001" => data <= "000000";
				when "001011100001011010" => data <= "000000";
				when "001011100001011011" => data <= "000000";
				when "001011100001011100" => data <= "000000";
				when "001011100001011101" => data <= "000000";
				when "001011100001011110" => data <= "000000";
				when "001011100001011111" => data <= "000000";
				when "001011100001100000" => data <= "000000";
				when "001011100001100001" => data <= "000000";
				when "001011100001100010" => data <= "000000";
				when "001011100001100011" => data <= "000000";
				when "001011100001100100" => data <= "000000";
				when "001011100001100101" => data <= "000000";
				when "001011100001100110" => data <= "000000";
				when "001011100001100111" => data <= "000000";
				when "001011100001101000" => data <= "000000";
				when "001011100001101001" => data <= "000000";
				when "001011100001101010" => data <= "000000";
				when "001011100001101011" => data <= "000000";
				when "001011100001101100" => data <= "000000";
				when "001011100001101101" => data <= "000000";
				when "001011100001101110" => data <= "000000";
				when "001011100001101111" => data <= "000000";
				when "001011100001110000" => data <= "000000";
				when "001011100001110001" => data <= "000000";
				when "001011100001110010" => data <= "000000";
				when "001011100001110011" => data <= "000000";
				when "001011100001110100" => data <= "000000";
				when "001011100001110101" => data <= "000000";
				when "001011100001110110" => data <= "000000";
				when "001011100001110111" => data <= "000000";
				when "001011100001111000" => data <= "000000";
				when "001011100001111001" => data <= "000000";
				when "001011100001111010" => data <= "000000";
				when "001011100001111011" => data <= "000000";
				when "001011100001111100" => data <= "000000";
				when "001011100001111101" => data <= "000000";
				when "001011100001111110" => data <= "000000";
				when "001011100001111111" => data <= "000000";
				when "001011100010000000" => data <= "000000";
				when "001011100010000001" => data <= "000000";
				when "001011100010000010" => data <= "000000";
				when "001011100010000011" => data <= "000000";
				when "001011100010000100" => data <= "000000";
				when "001011100010000101" => data <= "000000";
				when "001011100010000110" => data <= "000000";
				when "001011100010000111" => data <= "000000";
				when "001011100010001000" => data <= "000000";
				when "001011100010001001" => data <= "000000";
				when "001011100010001010" => data <= "000000";
				when "001011100010001011" => data <= "000000";
				when "001011100010001100" => data <= "000000";
				when "001011100010001101" => data <= "000000";
				when "001011100010001110" => data <= "000000";
				when "001011100010001111" => data <= "000000";
				when "001011100010010000" => data <= "000000";
				when "001011100010010001" => data <= "000000";
				when "001011100010010010" => data <= "000000";
				when "001011100010010011" => data <= "000000";
				when "001011100010010100" => data <= "000000";
				when "001011100010010101" => data <= "000000";
				when "001011100010010110" => data <= "000000";
				when "001011100010010111" => data <= "000000";
				when "001011100010011000" => data <= "000000";
				when "001011100010011001" => data <= "000000";
				when "001011100010011010" => data <= "000000";
				when "001011100010011011" => data <= "000000";
				when "001011100010011100" => data <= "000000";
				when "001011100010011101" => data <= "000000";
				when "001011100010011110" => data <= "000000";
				when "001011100010011111" => data <= "000000";
				when "001011101000000000" => data <= "000000";
				when "001011101000000001" => data <= "000000";
				when "001011101000000010" => data <= "000000";
				when "001011101000000011" => data <= "000000";
				when "001011101000000100" => data <= "000000";
				when "001011101000000101" => data <= "000000";
				when "001011101000000110" => data <= "000000";
				when "001011101000000111" => data <= "000000";
				when "001011101000001000" => data <= "000000";
				when "001011101000001001" => data <= "000000";
				when "001011101000001010" => data <= "000000";
				when "001011101000001011" => data <= "000000";
				when "001011101000001100" => data <= "000000";
				when "001011101000001101" => data <= "000000";
				when "001011101000001110" => data <= "000000";
				when "001011101000001111" => data <= "000000";
				when "001011101000010000" => data <= "000000";
				when "001011101000010001" => data <= "000000";
				when "001011101000010010" => data <= "000000";
				when "001011101000010011" => data <= "000000";
				when "001011101000010100" => data <= "000000";
				when "001011101000010101" => data <= "000000";
				when "001011101000010110" => data <= "000000";
				when "001011101000010111" => data <= "000000";
				when "001011101000011000" => data <= "000000";
				when "001011101000011001" => data <= "000000";
				when "001011101000011010" => data <= "000000";
				when "001011101000011011" => data <= "000000";
				when "001011101000011100" => data <= "000000";
				when "001011101000011101" => data <= "000000";
				when "001011101000011110" => data <= "000000";
				when "001011101000011111" => data <= "000000";
				when "001011101000100000" => data <= "000000";
				when "001011101000100001" => data <= "000000";
				when "001011101000100010" => data <= "000000";
				when "001011101000100011" => data <= "000000";
				when "001011101000100100" => data <= "000000";
				when "001011101000100101" => data <= "000000";
				when "001011101000100110" => data <= "000000";
				when "001011101000100111" => data <= "000000";
				when "001011101000101000" => data <= "000000";
				when "001011101000101001" => data <= "000000";
				when "001011101000101010" => data <= "000000";
				when "001011101000101011" => data <= "000000";
				when "001011101000101100" => data <= "000000";
				when "001011101000101101" => data <= "000000";
				when "001011101000101110" => data <= "000000";
				when "001011101000101111" => data <= "000000";
				when "001011101000110000" => data <= "000000";
				when "001011101000110001" => data <= "000000";
				when "001011101000110010" => data <= "000000";
				when "001011101000110011" => data <= "000000";
				when "001011101000110100" => data <= "000000";
				when "001011101000110101" => data <= "000000";
				when "001011101000110110" => data <= "000000";
				when "001011101000110111" => data <= "000000";
				when "001011101000111000" => data <= "000000";
				when "001011101000111001" => data <= "000000";
				when "001011101000111010" => data <= "000000";
				when "001011101000111011" => data <= "000000";
				when "001011101000111100" => data <= "000000";
				when "001011101000111101" => data <= "000000";
				when "001011101000111110" => data <= "000000";
				when "001011101000111111" => data <= "000000";
				when "001011101001000000" => data <= "000000";
				when "001011101001000001" => data <= "000000";
				when "001011101001000010" => data <= "000000";
				when "001011101001000011" => data <= "000000";
				when "001011101001000100" => data <= "000000";
				when "001011101001000101" => data <= "000000";
				when "001011101001000110" => data <= "000000";
				when "001011101001000111" => data <= "000000";
				when "001011101001001000" => data <= "000000";
				when "001011101001001001" => data <= "000000";
				when "001011101001001010" => data <= "000000";
				when "001011101001001011" => data <= "000000";
				when "001011101001001100" => data <= "000000";
				when "001011101001001101" => data <= "000000";
				when "001011101001001110" => data <= "000000";
				when "001011101001001111" => data <= "000000";
				when "001011101001010000" => data <= "000000";
				when "001011101001010001" => data <= "000000";
				when "001011101001010010" => data <= "000000";
				when "001011101001010011" => data <= "000000";
				when "001011101001010100" => data <= "000000";
				when "001011101001010101" => data <= "000000";
				when "001011101001010110" => data <= "000000";
				when "001011101001010111" => data <= "000000";
				when "001011101001011000" => data <= "000000";
				when "001011101001011001" => data <= "000000";
				when "001011101001011010" => data <= "000000";
				when "001011101001011011" => data <= "000000";
				when "001011101001011100" => data <= "000000";
				when "001011101001011101" => data <= "000000";
				when "001011101001011110" => data <= "000000";
				when "001011101001011111" => data <= "000000";
				when "001011101001100000" => data <= "000000";
				when "001011101001100001" => data <= "000000";
				when "001011101001100010" => data <= "000000";
				when "001011101001100011" => data <= "000000";
				when "001011101001100100" => data <= "000000";
				when "001011101001100101" => data <= "000000";
				when "001011101001100110" => data <= "000000";
				when "001011101001100111" => data <= "000000";
				when "001011101001101000" => data <= "000000";
				when "001011101001101001" => data <= "000000";
				when "001011101001101010" => data <= "000000";
				when "001011101001101011" => data <= "000000";
				when "001011101001101100" => data <= "000000";
				when "001011101001101101" => data <= "000000";
				when "001011101001101110" => data <= "000000";
				when "001011101001101111" => data <= "000000";
				when "001011101001110000" => data <= "000000";
				when "001011101001110001" => data <= "000000";
				when "001011101001110010" => data <= "000000";
				when "001011101001110011" => data <= "000000";
				when "001011101001110100" => data <= "000000";
				when "001011101001110101" => data <= "000000";
				when "001011101001110110" => data <= "000000";
				when "001011101001110111" => data <= "000000";
				when "001011101001111000" => data <= "000000";
				when "001011101001111001" => data <= "000000";
				when "001011101001111010" => data <= "000000";
				when "001011101001111011" => data <= "000000";
				when "001011101001111100" => data <= "000000";
				when "001011101001111101" => data <= "000000";
				when "001011101001111110" => data <= "000000";
				when "001011101001111111" => data <= "000000";
				when "001011101010000000" => data <= "000000";
				when "001011101010000001" => data <= "000000";
				when "001011101010000010" => data <= "000000";
				when "001011101010000011" => data <= "000000";
				when "001011101010000100" => data <= "000000";
				when "001011101010000101" => data <= "000000";
				when "001011101010000110" => data <= "000000";
				when "001011101010000111" => data <= "000000";
				when "001011101010001000" => data <= "000000";
				when "001011101010001001" => data <= "000000";
				when "001011101010001010" => data <= "000000";
				when "001011101010001011" => data <= "000000";
				when "001011101010001100" => data <= "000000";
				when "001011101010001101" => data <= "000000";
				when "001011101010001110" => data <= "000000";
				when "001011101010001111" => data <= "000000";
				when "001011101010010000" => data <= "000000";
				when "001011101010010001" => data <= "000000";
				when "001011101010010010" => data <= "000000";
				when "001011101010010011" => data <= "000000";
				when "001011101010010100" => data <= "000000";
				when "001011101010010101" => data <= "000000";
				when "001011101010010110" => data <= "000000";
				when "001011101010010111" => data <= "000000";
				when "001011101010011000" => data <= "000000";
				when "001011101010011001" => data <= "000000";
				when "001011101010011010" => data <= "000000";
				when "001011101010011011" => data <= "000000";
				when "001011101010011100" => data <= "000000";
				when "001011101010011101" => data <= "000000";
				when "001011101010011110" => data <= "000000";
				when "001011101010011111" => data <= "000000";
				when "001011110000000000" => data <= "000000";
				when "001011110000000001" => data <= "000000";
				when "001011110000000010" => data <= "000000";
				when "001011110000000011" => data <= "000000";
				when "001011110000000100" => data <= "000000";
				when "001011110000000101" => data <= "000000";
				when "001011110000000110" => data <= "000000";
				when "001011110000000111" => data <= "000000";
				when "001011110000001000" => data <= "000000";
				when "001011110000001001" => data <= "000000";
				when "001011110000001010" => data <= "000000";
				when "001011110000001011" => data <= "000000";
				when "001011110000001100" => data <= "000000";
				when "001011110000001101" => data <= "000000";
				when "001011110000001110" => data <= "000000";
				when "001011110000001111" => data <= "000000";
				when "001011110000010000" => data <= "000000";
				when "001011110000010001" => data <= "000000";
				when "001011110000010010" => data <= "000000";
				when "001011110000010011" => data <= "000000";
				when "001011110000010100" => data <= "000000";
				when "001011110000010101" => data <= "000000";
				when "001011110000010110" => data <= "000000";
				when "001011110000010111" => data <= "000000";
				when "001011110000011000" => data <= "000000";
				when "001011110000011001" => data <= "000000";
				when "001011110000011010" => data <= "000000";
				when "001011110000011011" => data <= "000000";
				when "001011110000011100" => data <= "000000";
				when "001011110000011101" => data <= "000000";
				when "001011110000011110" => data <= "000000";
				when "001011110000011111" => data <= "000000";
				when "001011110000100000" => data <= "000000";
				when "001011110000100001" => data <= "000000";
				when "001011110000100010" => data <= "000000";
				when "001011110000100011" => data <= "000000";
				when "001011110000100100" => data <= "000000";
				when "001011110000100101" => data <= "000000";
				when "001011110000100110" => data <= "000000";
				when "001011110000100111" => data <= "000000";
				when "001011110000101000" => data <= "000000";
				when "001011110000101001" => data <= "000000";
				when "001011110000101010" => data <= "000000";
				when "001011110000101011" => data <= "000000";
				when "001011110000101100" => data <= "000000";
				when "001011110000101101" => data <= "000000";
				when "001011110000101110" => data <= "000000";
				when "001011110000101111" => data <= "000000";
				when "001011110000110000" => data <= "000000";
				when "001011110000110001" => data <= "000000";
				when "001011110000110010" => data <= "000000";
				when "001011110000110011" => data <= "000000";
				when "001011110000110100" => data <= "000000";
				when "001011110000110101" => data <= "000000";
				when "001011110000110110" => data <= "000000";
				when "001011110000110111" => data <= "000000";
				when "001011110000111000" => data <= "000000";
				when "001011110000111001" => data <= "000000";
				when "001011110000111010" => data <= "000000";
				when "001011110000111011" => data <= "000000";
				when "001011110000111100" => data <= "000000";
				when "001011110000111101" => data <= "000000";
				when "001011110000111110" => data <= "000000";
				when "001011110000111111" => data <= "000000";
				when "001011110001000000" => data <= "000000";
				when "001011110001000001" => data <= "000000";
				when "001011110001000010" => data <= "000000";
				when "001011110001000011" => data <= "000000";
				when "001011110001000100" => data <= "000000";
				when "001011110001000101" => data <= "000000";
				when "001011110001000110" => data <= "000000";
				when "001011110001000111" => data <= "000000";
				when "001011110001001000" => data <= "000000";
				when "001011110001001001" => data <= "000000";
				when "001011110001001010" => data <= "000000";
				when "001011110001001011" => data <= "000000";
				when "001011110001001100" => data <= "000000";
				when "001011110001001101" => data <= "000000";
				when "001011110001001110" => data <= "000000";
				when "001011110001001111" => data <= "000000";
				when "001011110001010000" => data <= "000000";
				when "001011110001010001" => data <= "000000";
				when "001011110001010010" => data <= "000000";
				when "001011110001010011" => data <= "000000";
				when "001011110001010100" => data <= "000000";
				when "001011110001010101" => data <= "000000";
				when "001011110001010110" => data <= "000000";
				when "001011110001010111" => data <= "000000";
				when "001011110001011000" => data <= "000000";
				when "001011110001011001" => data <= "000000";
				when "001011110001011010" => data <= "000000";
				when "001011110001011011" => data <= "000000";
				when "001011110001011100" => data <= "000000";
				when "001011110001011101" => data <= "000000";
				when "001011110001011110" => data <= "000000";
				when "001011110001011111" => data <= "000000";
				when "001011110001100000" => data <= "000000";
				when "001011110001100001" => data <= "000000";
				when "001011110001100010" => data <= "000000";
				when "001011110001100011" => data <= "000000";
				when "001011110001100100" => data <= "000000";
				when "001011110001100101" => data <= "000000";
				when "001011110001100110" => data <= "000000";
				when "001011110001100111" => data <= "000000";
				when "001011110001101000" => data <= "000000";
				when "001011110001101001" => data <= "000000";
				when "001011110001101010" => data <= "000000";
				when "001011110001101011" => data <= "000000";
				when "001011110001101100" => data <= "000000";
				when "001011110001101101" => data <= "000000";
				when "001011110001101110" => data <= "000000";
				when "001011110001101111" => data <= "000000";
				when "001011110001110000" => data <= "000000";
				when "001011110001110001" => data <= "000000";
				when "001011110001110010" => data <= "000000";
				when "001011110001110011" => data <= "000000";
				when "001011110001110100" => data <= "000000";
				when "001011110001110101" => data <= "000000";
				when "001011110001110110" => data <= "000000";
				when "001011110001110111" => data <= "000000";
				when "001011110001111000" => data <= "000000";
				when "001011110001111001" => data <= "000000";
				when "001011110001111010" => data <= "000000";
				when "001011110001111011" => data <= "000000";
				when "001011110001111100" => data <= "000000";
				when "001011110001111101" => data <= "000000";
				when "001011110001111110" => data <= "000000";
				when "001011110001111111" => data <= "000000";
				when "001011110010000000" => data <= "000000";
				when "001011110010000001" => data <= "000000";
				when "001011110010000010" => data <= "000000";
				when "001011110010000011" => data <= "000000";
				when "001011110010000100" => data <= "000000";
				when "001011110010000101" => data <= "000000";
				when "001011110010000110" => data <= "000000";
				when "001011110010000111" => data <= "000000";
				when "001011110010001000" => data <= "000000";
				when "001011110010001001" => data <= "000000";
				when "001011110010001010" => data <= "000000";
				when "001011110010001011" => data <= "000000";
				when "001011110010001100" => data <= "000000";
				when "001011110010001101" => data <= "000000";
				when "001011110010001110" => data <= "000000";
				when "001011110010001111" => data <= "000000";
				when "001011110010010000" => data <= "000000";
				when "001011110010010001" => data <= "000000";
				when "001011110010010010" => data <= "000000";
				when "001011110010010011" => data <= "000000";
				when "001011110010010100" => data <= "000000";
				when "001011110010010101" => data <= "000000";
				when "001011110010010110" => data <= "000000";
				when "001011110010010111" => data <= "000000";
				when "001011110010011000" => data <= "000000";
				when "001011110010011001" => data <= "000000";
				when "001011110010011010" => data <= "000000";
				when "001011110010011011" => data <= "000000";
				when "001011110010011100" => data <= "000000";
				when "001011110010011101" => data <= "000000";
				when "001011110010011110" => data <= "000000";
				when "001011110010011111" => data <= "000000";
				when "001011111000000000" => data <= "000000";
				when "001011111000000001" => data <= "000000";
				when "001011111000000010" => data <= "000000";
				when "001011111000000011" => data <= "000000";
				when "001011111000000100" => data <= "000000";
				when "001011111000000101" => data <= "000000";
				when "001011111000000110" => data <= "000000";
				when "001011111000000111" => data <= "000000";
				when "001011111000001000" => data <= "000000";
				when "001011111000001001" => data <= "000000";
				when "001011111000001010" => data <= "000000";
				when "001011111000001011" => data <= "000000";
				when "001011111000001100" => data <= "000000";
				when "001011111000001101" => data <= "000000";
				when "001011111000001110" => data <= "000000";
				when "001011111000001111" => data <= "000000";
				when "001011111000010000" => data <= "000000";
				when "001011111000010001" => data <= "000000";
				when "001011111000010010" => data <= "000000";
				when "001011111000010011" => data <= "000000";
				when "001011111000010100" => data <= "000000";
				when "001011111000010101" => data <= "000000";
				when "001011111000010110" => data <= "000000";
				when "001011111000010111" => data <= "000000";
				when "001011111000011000" => data <= "000000";
				when "001011111000011001" => data <= "000000";
				when "001011111000011010" => data <= "000000";
				when "001011111000011011" => data <= "000000";
				when "001011111000011100" => data <= "000000";
				when "001011111000011101" => data <= "000000";
				when "001011111000011110" => data <= "000000";
				when "001011111000011111" => data <= "000000";
				when "001011111000100000" => data <= "000000";
				when "001011111000100001" => data <= "000000";
				when "001011111000100010" => data <= "000000";
				when "001011111000100011" => data <= "000000";
				when "001011111000100100" => data <= "000000";
				when "001011111000100101" => data <= "000000";
				when "001011111000100110" => data <= "000000";
				when "001011111000100111" => data <= "000000";
				when "001011111000101000" => data <= "000000";
				when "001011111000101001" => data <= "000000";
				when "001011111000101010" => data <= "000000";
				when "001011111000101011" => data <= "000000";
				when "001011111000101100" => data <= "000000";
				when "001011111000101101" => data <= "000000";
				when "001011111000101110" => data <= "000000";
				when "001011111000101111" => data <= "000000";
				when "001011111000110000" => data <= "000000";
				when "001011111000110001" => data <= "000000";
				when "001011111000110010" => data <= "000000";
				when "001011111000110011" => data <= "000000";
				when "001011111000110100" => data <= "000000";
				when "001011111000110101" => data <= "000000";
				when "001011111000110110" => data <= "000000";
				when "001011111000110111" => data <= "000000";
				when "001011111000111000" => data <= "000000";
				when "001011111000111001" => data <= "000000";
				when "001011111000111010" => data <= "000000";
				when "001011111000111011" => data <= "000000";
				when "001011111000111100" => data <= "000000";
				when "001011111000111101" => data <= "000000";
				when "001011111000111110" => data <= "000000";
				when "001011111000111111" => data <= "000000";
				when "001011111001000000" => data <= "000000";
				when "001011111001000001" => data <= "000000";
				when "001011111001000010" => data <= "000000";
				when "001011111001000011" => data <= "000000";
				when "001011111001000100" => data <= "000000";
				when "001011111001000101" => data <= "000000";
				when "001011111001000110" => data <= "000000";
				when "001011111001000111" => data <= "000000";
				when "001011111001001000" => data <= "000000";
				when "001011111001001001" => data <= "000000";
				when "001011111001001010" => data <= "000000";
				when "001011111001001011" => data <= "000000";
				when "001011111001001100" => data <= "000000";
				when "001011111001001101" => data <= "000000";
				when "001011111001001110" => data <= "000000";
				when "001011111001001111" => data <= "000000";
				when "001011111001010000" => data <= "000000";
				when "001011111001010001" => data <= "000000";
				when "001011111001010010" => data <= "000000";
				when "001011111001010011" => data <= "000000";
				when "001011111001010100" => data <= "000000";
				when "001011111001010101" => data <= "000000";
				when "001011111001010110" => data <= "000000";
				when "001011111001010111" => data <= "000000";
				when "001011111001011000" => data <= "000000";
				when "001011111001011001" => data <= "000000";
				when "001011111001011010" => data <= "000000";
				when "001011111001011011" => data <= "000000";
				when "001011111001011100" => data <= "000000";
				when "001011111001011101" => data <= "000000";
				when "001011111001011110" => data <= "000000";
				when "001011111001011111" => data <= "000000";
				when "001011111001100000" => data <= "000000";
				when "001011111001100001" => data <= "000000";
				when "001011111001100010" => data <= "000000";
				when "001011111001100011" => data <= "000000";
				when "001011111001100100" => data <= "000000";
				when "001011111001100101" => data <= "000000";
				when "001011111001100110" => data <= "000000";
				when "001011111001100111" => data <= "000000";
				when "001011111001101000" => data <= "000000";
				when "001011111001101001" => data <= "000000";
				when "001011111001101010" => data <= "000000";
				when "001011111001101011" => data <= "000000";
				when "001011111001101100" => data <= "000000";
				when "001011111001101101" => data <= "000000";
				when "001011111001101110" => data <= "000000";
				when "001011111001101111" => data <= "000000";
				when "001011111001110000" => data <= "000000";
				when "001011111001110001" => data <= "000000";
				when "001011111001110010" => data <= "000000";
				when "001011111001110011" => data <= "000000";
				when "001011111001110100" => data <= "000000";
				when "001011111001110101" => data <= "000000";
				when "001011111001110110" => data <= "000000";
				when "001011111001110111" => data <= "000000";
				when "001011111001111000" => data <= "000000";
				when "001011111001111001" => data <= "000000";
				when "001011111001111010" => data <= "000000";
				when "001011111001111011" => data <= "000000";
				when "001011111001111100" => data <= "000000";
				when "001011111001111101" => data <= "000000";
				when "001011111001111110" => data <= "000000";
				when "001011111001111111" => data <= "000000";
				when "001011111010000000" => data <= "000000";
				when "001011111010000001" => data <= "000000";
				when "001011111010000010" => data <= "000000";
				when "001011111010000011" => data <= "000000";
				when "001011111010000100" => data <= "000000";
				when "001011111010000101" => data <= "000000";
				when "001011111010000110" => data <= "000000";
				when "001011111010000111" => data <= "000000";
				when "001011111010001000" => data <= "000000";
				when "001011111010001001" => data <= "000000";
				when "001011111010001010" => data <= "000000";
				when "001011111010001011" => data <= "000000";
				when "001011111010001100" => data <= "000000";
				when "001011111010001101" => data <= "000000";
				when "001011111010001110" => data <= "000000";
				when "001011111010001111" => data <= "000000";
				when "001011111010010000" => data <= "000000";
				when "001011111010010001" => data <= "000000";
				when "001011111010010010" => data <= "000000";
				when "001011111010010011" => data <= "000000";
				when "001011111010010100" => data <= "000000";
				when "001011111010010101" => data <= "000000";
				when "001011111010010110" => data <= "000000";
				when "001011111010010111" => data <= "000000";
				when "001011111010011000" => data <= "000000";
				when "001011111010011001" => data <= "000000";
				when "001011111010011010" => data <= "000000";
				when "001011111010011011" => data <= "000000";
				when "001011111010011100" => data <= "000000";
				when "001011111010011101" => data <= "000000";
				when "001011111010011110" => data <= "000000";
				when "001011111010011111" => data <= "000000";
				when "001100000000000000" => data <= "000000";
				when "001100000000000001" => data <= "000000";
				when "001100000000000010" => data <= "000000";
				when "001100000000000011" => data <= "000000";
				when "001100000000000100" => data <= "000000";
				when "001100000000000101" => data <= "000000";
				when "001100000000000110" => data <= "000000";
				when "001100000000000111" => data <= "000000";
				when "001100000000001000" => data <= "000000";
				when "001100000000001001" => data <= "000000";
				when "001100000000001010" => data <= "000000";
				when "001100000000001011" => data <= "000000";
				when "001100000000001100" => data <= "000000";
				when "001100000000001101" => data <= "000000";
				when "001100000000001110" => data <= "000000";
				when "001100000000001111" => data <= "000000";
				when "001100000000010000" => data <= "000000";
				when "001100000000010001" => data <= "000000";
				when "001100000000010010" => data <= "000000";
				when "001100000000010011" => data <= "000000";
				when "001100000000010100" => data <= "000000";
				when "001100000000010101" => data <= "000000";
				when "001100000000010110" => data <= "000000";
				when "001100000000010111" => data <= "000000";
				when "001100000000011000" => data <= "000000";
				when "001100000000011001" => data <= "000000";
				when "001100000000011010" => data <= "000000";
				when "001100000000011011" => data <= "000000";
				when "001100000000011100" => data <= "000000";
				when "001100000000011101" => data <= "000000";
				when "001100000000011110" => data <= "000000";
				when "001100000000011111" => data <= "000000";
				when "001100000000100000" => data <= "000000";
				when "001100000000100001" => data <= "000000";
				when "001100000000100010" => data <= "000000";
				when "001100000000100011" => data <= "000000";
				when "001100000000100100" => data <= "000000";
				when "001100000000100101" => data <= "000000";
				when "001100000000100110" => data <= "000000";
				when "001100000000100111" => data <= "000000";
				when "001100000000101000" => data <= "000000";
				when "001100000000101001" => data <= "000000";
				when "001100000000101010" => data <= "000000";
				when "001100000000101011" => data <= "000000";
				when "001100000000101100" => data <= "000000";
				when "001100000000101101" => data <= "000000";
				when "001100000000101110" => data <= "000000";
				when "001100000000101111" => data <= "000000";
				when "001100000000110000" => data <= "000000";
				when "001100000000110001" => data <= "000000";
				when "001100000000110010" => data <= "000000";
				when "001100000000110011" => data <= "000000";
				when "001100000000110100" => data <= "000000";
				when "001100000000110101" => data <= "000000";
				when "001100000000110110" => data <= "000000";
				when "001100000000110111" => data <= "000000";
				when "001100000000111000" => data <= "000000";
				when "001100000000111001" => data <= "000000";
				when "001100000000111010" => data <= "000000";
				when "001100000000111011" => data <= "000000";
				when "001100000000111100" => data <= "000000";
				when "001100000000111101" => data <= "000000";
				when "001100000000111110" => data <= "000000";
				when "001100000000111111" => data <= "000000";
				when "001100000001000000" => data <= "000000";
				when "001100000001000001" => data <= "000000";
				when "001100000001000010" => data <= "000000";
				when "001100000001000011" => data <= "000000";
				when "001100000001000100" => data <= "000000";
				when "001100000001000101" => data <= "000000";
				when "001100000001000110" => data <= "000000";
				when "001100000001000111" => data <= "000000";
				when "001100000001001000" => data <= "000000";
				when "001100000001001001" => data <= "000000";
				when "001100000001001010" => data <= "000000";
				when "001100000001001011" => data <= "000000";
				when "001100000001001100" => data <= "000000";
				when "001100000001001101" => data <= "000000";
				when "001100000001001110" => data <= "000000";
				when "001100000001001111" => data <= "000000";
				when "001100000001010000" => data <= "000000";
				when "001100000001010001" => data <= "000000";
				when "001100000001010010" => data <= "000000";
				when "001100000001010011" => data <= "000000";
				when "001100000001010100" => data <= "000000";
				when "001100000001010101" => data <= "000000";
				when "001100000001010110" => data <= "000000";
				when "001100000001010111" => data <= "000000";
				when "001100000001011000" => data <= "000000";
				when "001100000001011001" => data <= "000000";
				when "001100000001011010" => data <= "000000";
				when "001100000001011011" => data <= "000000";
				when "001100000001011100" => data <= "000000";
				when "001100000001011101" => data <= "000000";
				when "001100000001011110" => data <= "000000";
				when "001100000001011111" => data <= "000000";
				when "001100000001100000" => data <= "000000";
				when "001100000001100001" => data <= "000000";
				when "001100000001100010" => data <= "000000";
				when "001100000001100011" => data <= "000000";
				when "001100000001100100" => data <= "000000";
				when "001100000001100101" => data <= "000000";
				when "001100000001100110" => data <= "000000";
				when "001100000001100111" => data <= "000000";
				when "001100000001101000" => data <= "000000";
				when "001100000001101001" => data <= "000000";
				when "001100000001101010" => data <= "000000";
				when "001100000001101011" => data <= "000000";
				when "001100000001101100" => data <= "000000";
				when "001100000001101101" => data <= "000000";
				when "001100000001101110" => data <= "000000";
				when "001100000001101111" => data <= "000000";
				when "001100000001110000" => data <= "000000";
				when "001100000001110001" => data <= "000000";
				when "001100000001110010" => data <= "000000";
				when "001100000001110011" => data <= "000000";
				when "001100000001110100" => data <= "000000";
				when "001100000001110101" => data <= "000000";
				when "001100000001110110" => data <= "000000";
				when "001100000001110111" => data <= "000000";
				when "001100000001111000" => data <= "000000";
				when "001100000001111001" => data <= "000000";
				when "001100000001111010" => data <= "000000";
				when "001100000001111011" => data <= "000000";
				when "001100000001111100" => data <= "000000";
				when "001100000001111101" => data <= "000000";
				when "001100000001111110" => data <= "000000";
				when "001100000001111111" => data <= "000000";
				when "001100000010000000" => data <= "000000";
				when "001100000010000001" => data <= "000000";
				when "001100000010000010" => data <= "000000";
				when "001100000010000011" => data <= "000000";
				when "001100000010000100" => data <= "000000";
				when "001100000010000101" => data <= "000000";
				when "001100000010000110" => data <= "000000";
				when "001100000010000111" => data <= "000000";
				when "001100000010001000" => data <= "000000";
				when "001100000010001001" => data <= "000000";
				when "001100000010001010" => data <= "000000";
				when "001100000010001011" => data <= "000000";
				when "001100000010001100" => data <= "000000";
				when "001100000010001101" => data <= "000000";
				when "001100000010001110" => data <= "000000";
				when "001100000010001111" => data <= "000000";
				when "001100000010010000" => data <= "000000";
				when "001100000010010001" => data <= "000000";
				when "001100000010010010" => data <= "000000";
				when "001100000010010011" => data <= "000000";
				when "001100000010010100" => data <= "000000";
				when "001100000010010101" => data <= "000000";
				when "001100000010010110" => data <= "000000";
				when "001100000010010111" => data <= "000000";
				when "001100000010011000" => data <= "000000";
				when "001100000010011001" => data <= "000000";
				when "001100000010011010" => data <= "000000";
				when "001100000010011011" => data <= "000000";
				when "001100000010011100" => data <= "000000";
				when "001100000010011101" => data <= "000000";
				when "001100000010011110" => data <= "000000";
				when "001100000010011111" => data <= "000000";
				when "001100001000000000" => data <= "000000";
				when "001100001000000001" => data <= "000000";
				when "001100001000000010" => data <= "000000";
				when "001100001000000011" => data <= "000000";
				when "001100001000000100" => data <= "000000";
				when "001100001000000101" => data <= "000000";
				when "001100001000000110" => data <= "000000";
				when "001100001000000111" => data <= "000000";
				when "001100001000001000" => data <= "000000";
				when "001100001000001001" => data <= "000000";
				when "001100001000001010" => data <= "000000";
				when "001100001000001011" => data <= "000000";
				when "001100001000001100" => data <= "000000";
				when "001100001000001101" => data <= "000000";
				when "001100001000001110" => data <= "000000";
				when "001100001000001111" => data <= "000000";
				when "001100001000010000" => data <= "000000";
				when "001100001000010001" => data <= "000000";
				when "001100001000010010" => data <= "000000";
				when "001100001000010011" => data <= "000000";
				when "001100001000010100" => data <= "000000";
				when "001100001000010101" => data <= "000000";
				when "001100001000010110" => data <= "000000";
				when "001100001000010111" => data <= "000000";
				when "001100001000011000" => data <= "000000";
				when "001100001000011001" => data <= "000000";
				when "001100001000011010" => data <= "000000";
				when "001100001000011011" => data <= "000000";
				when "001100001000011100" => data <= "000000";
				when "001100001000011101" => data <= "000000";
				when "001100001000011110" => data <= "000000";
				when "001100001000011111" => data <= "000000";
				when "001100001000100000" => data <= "000000";
				when "001100001000100001" => data <= "000000";
				when "001100001000100010" => data <= "000000";
				when "001100001000100011" => data <= "000000";
				when "001100001000100100" => data <= "000000";
				when "001100001000100101" => data <= "000000";
				when "001100001000100110" => data <= "000000";
				when "001100001000100111" => data <= "000000";
				when "001100001000101000" => data <= "000000";
				when "001100001000101001" => data <= "000000";
				when "001100001000101010" => data <= "000000";
				when "001100001000101011" => data <= "000000";
				when "001100001000101100" => data <= "000000";
				when "001100001000101101" => data <= "000000";
				when "001100001000101110" => data <= "000000";
				when "001100001000101111" => data <= "000000";
				when "001100001000110000" => data <= "000000";
				when "001100001000110001" => data <= "000000";
				when "001100001000110010" => data <= "000000";
				when "001100001000110011" => data <= "000000";
				when "001100001000110100" => data <= "000000";
				when "001100001000110101" => data <= "000000";
				when "001100001000110110" => data <= "000000";
				when "001100001000110111" => data <= "000000";
				when "001100001000111000" => data <= "000000";
				when "001100001000111001" => data <= "000000";
				when "001100001000111010" => data <= "000000";
				when "001100001000111011" => data <= "000000";
				when "001100001000111100" => data <= "000000";
				when "001100001000111101" => data <= "000000";
				when "001100001000111110" => data <= "000000";
				when "001100001000111111" => data <= "000000";
				when "001100001001000000" => data <= "000000";
				when "001100001001000001" => data <= "000000";
				when "001100001001000010" => data <= "000000";
				when "001100001001000011" => data <= "000000";
				when "001100001001000100" => data <= "000000";
				when "001100001001000101" => data <= "000000";
				when "001100001001000110" => data <= "000000";
				when "001100001001000111" => data <= "000000";
				when "001100001001001000" => data <= "000000";
				when "001100001001001001" => data <= "000000";
				when "001100001001001010" => data <= "000000";
				when "001100001001001011" => data <= "000000";
				when "001100001001001100" => data <= "000000";
				when "001100001001001101" => data <= "000000";
				when "001100001001001110" => data <= "000000";
				when "001100001001001111" => data <= "000000";
				when "001100001001010000" => data <= "000000";
				when "001100001001010001" => data <= "000000";
				when "001100001001010010" => data <= "000000";
				when "001100001001010011" => data <= "000000";
				when "001100001001010100" => data <= "000000";
				when "001100001001010101" => data <= "000000";
				when "001100001001010110" => data <= "000000";
				when "001100001001010111" => data <= "000000";
				when "001100001001011000" => data <= "000000";
				when "001100001001011001" => data <= "000000";
				when "001100001001011010" => data <= "000000";
				when "001100001001011011" => data <= "000000";
				when "001100001001011100" => data <= "000000";
				when "001100001001011101" => data <= "000000";
				when "001100001001011110" => data <= "000000";
				when "001100001001011111" => data <= "000000";
				when "001100001001100000" => data <= "000000";
				when "001100001001100001" => data <= "000000";
				when "001100001001100010" => data <= "000000";
				when "001100001001100011" => data <= "000000";
				when "001100001001100100" => data <= "000000";
				when "001100001001100101" => data <= "000000";
				when "001100001001100110" => data <= "000000";
				when "001100001001100111" => data <= "000000";
				when "001100001001101000" => data <= "000000";
				when "001100001001101001" => data <= "000000";
				when "001100001001101010" => data <= "000000";
				when "001100001001101011" => data <= "000000";
				when "001100001001101100" => data <= "000000";
				when "001100001001101101" => data <= "000000";
				when "001100001001101110" => data <= "000000";
				when "001100001001101111" => data <= "000000";
				when "001100001001110000" => data <= "000000";
				when "001100001001110001" => data <= "000000";
				when "001100001001110010" => data <= "000000";
				when "001100001001110011" => data <= "000000";
				when "001100001001110100" => data <= "000000";
				when "001100001001110101" => data <= "000000";
				when "001100001001110110" => data <= "000000";
				when "001100001001110111" => data <= "000000";
				when "001100001001111000" => data <= "000000";
				when "001100001001111001" => data <= "000000";
				when "001100001001111010" => data <= "000000";
				when "001100001001111011" => data <= "000000";
				when "001100001001111100" => data <= "000000";
				when "001100001001111101" => data <= "000000";
				when "001100001001111110" => data <= "000000";
				when "001100001001111111" => data <= "000000";
				when "001100001010000000" => data <= "000000";
				when "001100001010000001" => data <= "000000";
				when "001100001010000010" => data <= "000000";
				when "001100001010000011" => data <= "000000";
				when "001100001010000100" => data <= "000000";
				when "001100001010000101" => data <= "000000";
				when "001100001010000110" => data <= "000000";
				when "001100001010000111" => data <= "000000";
				when "001100001010001000" => data <= "000000";
				when "001100001010001001" => data <= "000000";
				when "001100001010001010" => data <= "000000";
				when "001100001010001011" => data <= "000000";
				when "001100001010001100" => data <= "000000";
				when "001100001010001101" => data <= "000000";
				when "001100001010001110" => data <= "000000";
				when "001100001010001111" => data <= "000000";
				when "001100001010010000" => data <= "000000";
				when "001100001010010001" => data <= "000000";
				when "001100001010010010" => data <= "000000";
				when "001100001010010011" => data <= "000000";
				when "001100001010010100" => data <= "000000";
				when "001100001010010101" => data <= "000000";
				when "001100001010010110" => data <= "000000";
				when "001100001010010111" => data <= "000000";
				when "001100001010011000" => data <= "000000";
				when "001100001010011001" => data <= "000000";
				when "001100001010011010" => data <= "000000";
				when "001100001010011011" => data <= "000000";
				when "001100001010011100" => data <= "000000";
				when "001100001010011101" => data <= "000000";
				when "001100001010011110" => data <= "000000";
				when "001100001010011111" => data <= "000000";
				when "001100010000000000" => data <= "000000";
				when "001100010000000001" => data <= "000000";
				when "001100010000000010" => data <= "000000";
				when "001100010000000011" => data <= "000000";
				when "001100010000000100" => data <= "000000";
				when "001100010000000101" => data <= "000000";
				when "001100010000000110" => data <= "000000";
				when "001100010000000111" => data <= "000000";
				when "001100010000001000" => data <= "000000";
				when "001100010000001001" => data <= "000000";
				when "001100010000001010" => data <= "000000";
				when "001100010000001011" => data <= "000000";
				when "001100010000001100" => data <= "000000";
				when "001100010000001101" => data <= "000000";
				when "001100010000001110" => data <= "000000";
				when "001100010000001111" => data <= "000000";
				when "001100010000010000" => data <= "000000";
				when "001100010000010001" => data <= "000000";
				when "001100010000010010" => data <= "000000";
				when "001100010000010011" => data <= "000000";
				when "001100010000010100" => data <= "000000";
				when "001100010000010101" => data <= "000000";
				when "001100010000010110" => data <= "000000";
				when "001100010000010111" => data <= "000000";
				when "001100010000011000" => data <= "000000";
				when "001100010000011001" => data <= "000000";
				when "001100010000011010" => data <= "000000";
				when "001100010000011011" => data <= "000000";
				when "001100010000011100" => data <= "000000";
				when "001100010000011101" => data <= "000000";
				when "001100010000011110" => data <= "000000";
				when "001100010000011111" => data <= "000000";
				when "001100010000100000" => data <= "000000";
				when "001100010000100001" => data <= "000000";
				when "001100010000100010" => data <= "000000";
				when "001100010000100011" => data <= "000000";
				when "001100010000100100" => data <= "000000";
				when "001100010000100101" => data <= "000000";
				when "001100010000100110" => data <= "000000";
				when "001100010000100111" => data <= "000000";
				when "001100010000101000" => data <= "000000";
				when "001100010000101001" => data <= "000000";
				when "001100010000101010" => data <= "000000";
				when "001100010000101011" => data <= "000000";
				when "001100010000101100" => data <= "000000";
				when "001100010000101101" => data <= "000000";
				when "001100010000101110" => data <= "000000";
				when "001100010000101111" => data <= "000000";
				when "001100010000110000" => data <= "000000";
				when "001100010000110001" => data <= "000000";
				when "001100010000110010" => data <= "000000";
				when "001100010000110011" => data <= "000000";
				when "001100010000110100" => data <= "000000";
				when "001100010000110101" => data <= "000000";
				when "001100010000110110" => data <= "000000";
				when "001100010000110111" => data <= "000000";
				when "001100010000111000" => data <= "000000";
				when "001100010000111001" => data <= "000000";
				when "001100010000111010" => data <= "000000";
				when "001100010000111011" => data <= "000000";
				when "001100010000111100" => data <= "000000";
				when "001100010000111101" => data <= "000000";
				when "001100010000111110" => data <= "000000";
				when "001100010000111111" => data <= "000000";
				when "001100010001000000" => data <= "000000";
				when "001100010001000001" => data <= "000000";
				when "001100010001000010" => data <= "000000";
				when "001100010001000011" => data <= "000000";
				when "001100010001000100" => data <= "000000";
				when "001100010001000101" => data <= "000000";
				when "001100010001000110" => data <= "000000";
				when "001100010001000111" => data <= "000000";
				when "001100010001001000" => data <= "000000";
				when "001100010001001001" => data <= "000000";
				when "001100010001001010" => data <= "000000";
				when "001100010001001011" => data <= "000000";
				when "001100010001001100" => data <= "000000";
				when "001100010001001101" => data <= "000000";
				when "001100010001001110" => data <= "000000";
				when "001100010001001111" => data <= "000000";
				when "001100010001010000" => data <= "000000";
				when "001100010001010001" => data <= "000000";
				when "001100010001010010" => data <= "000000";
				when "001100010001010011" => data <= "000000";
				when "001100010001010100" => data <= "000000";
				when "001100010001010101" => data <= "000000";
				when "001100010001010110" => data <= "000000";
				when "001100010001010111" => data <= "000000";
				when "001100010001011000" => data <= "000000";
				when "001100010001011001" => data <= "000000";
				when "001100010001011010" => data <= "000000";
				when "001100010001011011" => data <= "000000";
				when "001100010001011100" => data <= "000000";
				when "001100010001011101" => data <= "000000";
				when "001100010001011110" => data <= "000000";
				when "001100010001011111" => data <= "000000";
				when "001100010001100000" => data <= "000000";
				when "001100010001100001" => data <= "000000";
				when "001100010001100010" => data <= "000000";
				when "001100010001100011" => data <= "000000";
				when "001100010001100100" => data <= "000000";
				when "001100010001100101" => data <= "000000";
				when "001100010001100110" => data <= "000000";
				when "001100010001100111" => data <= "000000";
				when "001100010001101000" => data <= "000000";
				when "001100010001101001" => data <= "000000";
				when "001100010001101010" => data <= "000000";
				when "001100010001101011" => data <= "000000";
				when "001100010001101100" => data <= "000000";
				when "001100010001101101" => data <= "000000";
				when "001100010001101110" => data <= "000000";
				when "001100010001101111" => data <= "000000";
				when "001100010001110000" => data <= "000000";
				when "001100010001110001" => data <= "000000";
				when "001100010001110010" => data <= "000000";
				when "001100010001110011" => data <= "000000";
				when "001100010001110100" => data <= "000000";
				when "001100010001110101" => data <= "000000";
				when "001100010001110110" => data <= "000000";
				when "001100010001110111" => data <= "000000";
				when "001100010001111000" => data <= "000000";
				when "001100010001111001" => data <= "000000";
				when "001100010001111010" => data <= "000000";
				when "001100010001111011" => data <= "000000";
				when "001100010001111100" => data <= "000000";
				when "001100010001111101" => data <= "000000";
				when "001100010001111110" => data <= "000000";
				when "001100010001111111" => data <= "000000";
				when "001100010010000000" => data <= "000000";
				when "001100010010000001" => data <= "000000";
				when "001100010010000010" => data <= "000000";
				when "001100010010000011" => data <= "000000";
				when "001100010010000100" => data <= "000000";
				when "001100010010000101" => data <= "000000";
				when "001100010010000110" => data <= "000000";
				when "001100010010000111" => data <= "000000";
				when "001100010010001000" => data <= "000000";
				when "001100010010001001" => data <= "000000";
				when "001100010010001010" => data <= "000000";
				when "001100010010001011" => data <= "000000";
				when "001100010010001100" => data <= "000000";
				when "001100010010001101" => data <= "000000";
				when "001100010010001110" => data <= "000000";
				when "001100010010001111" => data <= "000000";
				when "001100010010010000" => data <= "000000";
				when "001100010010010001" => data <= "000000";
				when "001100010010010010" => data <= "000000";
				when "001100010010010011" => data <= "000000";
				when "001100010010010100" => data <= "000000";
				when "001100010010010101" => data <= "000000";
				when "001100010010010110" => data <= "000000";
				when "001100010010010111" => data <= "000000";
				when "001100010010011000" => data <= "000000";
				when "001100010010011001" => data <= "000000";
				when "001100010010011010" => data <= "000000";
				when "001100010010011011" => data <= "000000";
				when "001100010010011100" => data <= "000000";
				when "001100010010011101" => data <= "000000";
				when "001100010010011110" => data <= "000000";
				when "001100010010011111" => data <= "000000";
				when "001100011000000000" => data <= "000000";
				when "001100011000000001" => data <= "000000";
				when "001100011000000010" => data <= "000000";
				when "001100011000000011" => data <= "000000";
				when "001100011000000100" => data <= "000000";
				when "001100011000000101" => data <= "000000";
				when "001100011000000110" => data <= "000000";
				when "001100011000000111" => data <= "000000";
				when "001100011000001000" => data <= "000000";
				when "001100011000001001" => data <= "000000";
				when "001100011000001010" => data <= "000000";
				when "001100011000001011" => data <= "000000";
				when "001100011000001100" => data <= "000000";
				when "001100011000001101" => data <= "000000";
				when "001100011000001110" => data <= "000000";
				when "001100011000001111" => data <= "000000";
				when "001100011000010000" => data <= "000000";
				when "001100011000010001" => data <= "000000";
				when "001100011000010010" => data <= "000000";
				when "001100011000010011" => data <= "000000";
				when "001100011000010100" => data <= "000000";
				when "001100011000010101" => data <= "000000";
				when "001100011000010110" => data <= "000000";
				when "001100011000010111" => data <= "000000";
				when "001100011000011000" => data <= "000000";
				when "001100011000011001" => data <= "000000";
				when "001100011000011010" => data <= "000000";
				when "001100011000011011" => data <= "000000";
				when "001100011000011100" => data <= "000000";
				when "001100011000011101" => data <= "000000";
				when "001100011000011110" => data <= "000000";
				when "001100011000011111" => data <= "000000";
				when "001100011000100000" => data <= "000000";
				when "001100011000100001" => data <= "000000";
				when "001100011000100010" => data <= "000000";
				when "001100011000100011" => data <= "000000";
				when "001100011000100100" => data <= "000000";
				when "001100011000100101" => data <= "000000";
				when "001100011000100110" => data <= "000000";
				when "001100011000100111" => data <= "000000";
				when "001100011000101000" => data <= "000000";
				when "001100011000101001" => data <= "000000";
				when "001100011000101010" => data <= "000000";
				when "001100011000101011" => data <= "000000";
				when "001100011000101100" => data <= "000000";
				when "001100011000101101" => data <= "000000";
				when "001100011000101110" => data <= "000000";
				when "001100011000101111" => data <= "000000";
				when "001100011000110000" => data <= "000000";
				when "001100011000110001" => data <= "000000";
				when "001100011000110010" => data <= "000000";
				when "001100011000110011" => data <= "000000";
				when "001100011000110100" => data <= "000000";
				when "001100011000110101" => data <= "000000";
				when "001100011000110110" => data <= "000000";
				when "001100011000110111" => data <= "000000";
				when "001100011000111000" => data <= "000000";
				when "001100011000111001" => data <= "000000";
				when "001100011000111010" => data <= "000000";
				when "001100011000111011" => data <= "000000";
				when "001100011000111100" => data <= "000000";
				when "001100011000111101" => data <= "000000";
				when "001100011000111110" => data <= "000000";
				when "001100011000111111" => data <= "000000";
				when "001100011001000000" => data <= "000000";
				when "001100011001000001" => data <= "000000";
				when "001100011001000010" => data <= "000000";
				when "001100011001000011" => data <= "000000";
				when "001100011001000100" => data <= "000000";
				when "001100011001000101" => data <= "000000";
				when "001100011001000110" => data <= "000000";
				when "001100011001000111" => data <= "000000";
				when "001100011001001000" => data <= "000000";
				when "001100011001001001" => data <= "000000";
				when "001100011001001010" => data <= "000000";
				when "001100011001001011" => data <= "000000";
				when "001100011001001100" => data <= "000000";
				when "001100011001001101" => data <= "000000";
				when "001100011001001110" => data <= "000000";
				when "001100011001001111" => data <= "000000";
				when "001100011001010000" => data <= "000000";
				when "001100011001010001" => data <= "000000";
				when "001100011001010010" => data <= "000000";
				when "001100011001010011" => data <= "000000";
				when "001100011001010100" => data <= "000000";
				when "001100011001010101" => data <= "000000";
				when "001100011001010110" => data <= "000000";
				when "001100011001010111" => data <= "000000";
				when "001100011001011000" => data <= "000000";
				when "001100011001011001" => data <= "000000";
				when "001100011001011010" => data <= "000000";
				when "001100011001011011" => data <= "000000";
				when "001100011001011100" => data <= "000000";
				when "001100011001011101" => data <= "000000";
				when "001100011001011110" => data <= "000000";
				when "001100011001011111" => data <= "000000";
				when "001100011001100000" => data <= "000000";
				when "001100011001100001" => data <= "000000";
				when "001100011001100010" => data <= "000000";
				when "001100011001100011" => data <= "000000";
				when "001100011001100100" => data <= "000000";
				when "001100011001100101" => data <= "000000";
				when "001100011001100110" => data <= "000000";
				when "001100011001100111" => data <= "000000";
				when "001100011001101000" => data <= "000000";
				when "001100011001101001" => data <= "000000";
				when "001100011001101010" => data <= "000000";
				when "001100011001101011" => data <= "000000";
				when "001100011001101100" => data <= "000000";
				when "001100011001101101" => data <= "000000";
				when "001100011001101110" => data <= "000000";
				when "001100011001101111" => data <= "000000";
				when "001100011001110000" => data <= "000000";
				when "001100011001110001" => data <= "000000";
				when "001100011001110010" => data <= "000000";
				when "001100011001110011" => data <= "000000";
				when "001100011001110100" => data <= "000000";
				when "001100011001110101" => data <= "000000";
				when "001100011001110110" => data <= "000000";
				when "001100011001110111" => data <= "000000";
				when "001100011001111000" => data <= "000000";
				when "001100011001111001" => data <= "000000";
				when "001100011001111010" => data <= "000000";
				when "001100011001111011" => data <= "000000";
				when "001100011001111100" => data <= "000000";
				when "001100011001111101" => data <= "000000";
				when "001100011001111110" => data <= "000000";
				when "001100011001111111" => data <= "000000";
				when "001100011010000000" => data <= "000000";
				when "001100011010000001" => data <= "000000";
				when "001100011010000010" => data <= "000000";
				when "001100011010000011" => data <= "000000";
				when "001100011010000100" => data <= "000000";
				when "001100011010000101" => data <= "000000";
				when "001100011010000110" => data <= "000000";
				when "001100011010000111" => data <= "000000";
				when "001100011010001000" => data <= "000000";
				when "001100011010001001" => data <= "000000";
				when "001100011010001010" => data <= "000000";
				when "001100011010001011" => data <= "000000";
				when "001100011010001100" => data <= "000000";
				when "001100011010001101" => data <= "000000";
				when "001100011010001110" => data <= "000000";
				when "001100011010001111" => data <= "000000";
				when "001100011010010000" => data <= "000000";
				when "001100011010010001" => data <= "000000";
				when "001100011010010010" => data <= "000000";
				when "001100011010010011" => data <= "000000";
				when "001100011010010100" => data <= "000000";
				when "001100011010010101" => data <= "000000";
				when "001100011010010110" => data <= "000000";
				when "001100011010010111" => data <= "000000";
				when "001100011010011000" => data <= "000000";
				when "001100011010011001" => data <= "000000";
				when "001100011010011010" => data <= "000000";
				when "001100011010011011" => data <= "000000";
				when "001100011010011100" => data <= "000000";
				when "001100011010011101" => data <= "000000";
				when "001100011010011110" => data <= "000000";
				when "001100011010011111" => data <= "000000";
				when "001100100000000000" => data <= "000000";
				when "001100100000000001" => data <= "000000";
				when "001100100000000010" => data <= "000000";
				when "001100100000000011" => data <= "000000";
				when "001100100000000100" => data <= "000000";
				when "001100100000000101" => data <= "000000";
				when "001100100000000110" => data <= "000000";
				when "001100100000000111" => data <= "000000";
				when "001100100000001000" => data <= "000000";
				when "001100100000001001" => data <= "000000";
				when "001100100000001010" => data <= "000000";
				when "001100100000001011" => data <= "000000";
				when "001100100000001100" => data <= "000000";
				when "001100100000001101" => data <= "000000";
				when "001100100000001110" => data <= "000000";
				when "001100100000001111" => data <= "000000";
				when "001100100000010000" => data <= "000000";
				when "001100100000010001" => data <= "000000";
				when "001100100000010010" => data <= "000000";
				when "001100100000010011" => data <= "000000";
				when "001100100000010100" => data <= "000000";
				when "001100100000010101" => data <= "000000";
				when "001100100000010110" => data <= "000000";
				when "001100100000010111" => data <= "000000";
				when "001100100000011000" => data <= "000000";
				when "001100100000011001" => data <= "000000";
				when "001100100000011010" => data <= "000000";
				when "001100100000011011" => data <= "000000";
				when "001100100000011100" => data <= "000000";
				when "001100100000011101" => data <= "000000";
				when "001100100000011110" => data <= "000000";
				when "001100100000011111" => data <= "000000";
				when "001100100000100000" => data <= "000000";
				when "001100100000100001" => data <= "000000";
				when "001100100000100010" => data <= "000000";
				when "001100100000100011" => data <= "000000";
				when "001100100000100100" => data <= "000000";
				when "001100100000100101" => data <= "000000";
				when "001100100000100110" => data <= "000000";
				when "001100100000100111" => data <= "000000";
				when "001100100000101000" => data <= "000000";
				when "001100100000101001" => data <= "000000";
				when "001100100000101010" => data <= "000000";
				when "001100100000101011" => data <= "000000";
				when "001100100000101100" => data <= "000000";
				when "001100100000101101" => data <= "000000";
				when "001100100000101110" => data <= "000000";
				when "001100100000101111" => data <= "000000";
				when "001100100000110000" => data <= "000000";
				when "001100100000110001" => data <= "000000";
				when "001100100000110010" => data <= "000000";
				when "001100100000110011" => data <= "000000";
				when "001100100000110100" => data <= "000000";
				when "001100100000110101" => data <= "000000";
				when "001100100000110110" => data <= "000000";
				when "001100100000110111" => data <= "000000";
				when "001100100000111000" => data <= "000000";
				when "001100100000111001" => data <= "000000";
				when "001100100000111010" => data <= "000000";
				when "001100100000111011" => data <= "000000";
				when "001100100000111100" => data <= "000000";
				when "001100100000111101" => data <= "000000";
				when "001100100000111110" => data <= "000000";
				when "001100100000111111" => data <= "000000";
				when "001100100001000000" => data <= "000000";
				when "001100100001000001" => data <= "000000";
				when "001100100001000010" => data <= "000000";
				when "001100100001000011" => data <= "000000";
				when "001100100001000100" => data <= "000000";
				when "001100100001000101" => data <= "000000";
				when "001100100001000110" => data <= "000000";
				when "001100100001000111" => data <= "000000";
				when "001100100001001000" => data <= "000000";
				when "001100100001001001" => data <= "000000";
				when "001100100001001010" => data <= "000000";
				when "001100100001001011" => data <= "000000";
				when "001100100001001100" => data <= "000000";
				when "001100100001001101" => data <= "000000";
				when "001100100001001110" => data <= "000000";
				when "001100100001001111" => data <= "000000";
				when "001100100001010000" => data <= "000000";
				when "001100100001010001" => data <= "000000";
				when "001100100001010010" => data <= "000000";
				when "001100100001010011" => data <= "000000";
				when "001100100001010100" => data <= "000000";
				when "001100100001010101" => data <= "000000";
				when "001100100001010110" => data <= "000000";
				when "001100100001010111" => data <= "000000";
				when "001100100001011000" => data <= "000000";
				when "001100100001011001" => data <= "000000";
				when "001100100001011010" => data <= "000000";
				when "001100100001011011" => data <= "000000";
				when "001100100001011100" => data <= "000000";
				when "001100100001011101" => data <= "000000";
				when "001100100001011110" => data <= "000000";
				when "001100100001011111" => data <= "000000";
				when "001100100001100000" => data <= "000000";
				when "001100100001100001" => data <= "000000";
				when "001100100001100010" => data <= "000000";
				when "001100100001100011" => data <= "000000";
				when "001100100001100100" => data <= "000000";
				when "001100100001100101" => data <= "000000";
				when "001100100001100110" => data <= "000000";
				when "001100100001100111" => data <= "000000";
				when "001100100001101000" => data <= "000000";
				when "001100100001101001" => data <= "000000";
				when "001100100001101010" => data <= "000000";
				when "001100100001101011" => data <= "000000";
				when "001100100001101100" => data <= "000000";
				when "001100100001101101" => data <= "000000";
				when "001100100001101110" => data <= "000000";
				when "001100100001101111" => data <= "000000";
				when "001100100001110000" => data <= "000000";
				when "001100100001110001" => data <= "000000";
				when "001100100001110010" => data <= "000000";
				when "001100100001110011" => data <= "000000";
				when "001100100001110100" => data <= "000000";
				when "001100100001110101" => data <= "000000";
				when "001100100001110110" => data <= "000000";
				when "001100100001110111" => data <= "000000";
				when "001100100001111000" => data <= "000000";
				when "001100100001111001" => data <= "000000";
				when "001100100001111010" => data <= "000000";
				when "001100100001111011" => data <= "000000";
				when "001100100001111100" => data <= "000000";
				when "001100100001111101" => data <= "000000";
				when "001100100001111110" => data <= "000000";
				when "001100100001111111" => data <= "000000";
				when "001100100010000000" => data <= "000000";
				when "001100100010000001" => data <= "000000";
				when "001100100010000010" => data <= "000000";
				when "001100100010000011" => data <= "000000";
				when "001100100010000100" => data <= "000000";
				when "001100100010000101" => data <= "000000";
				when "001100100010000110" => data <= "000000";
				when "001100100010000111" => data <= "000000";
				when "001100100010001000" => data <= "000000";
				when "001100100010001001" => data <= "000000";
				when "001100100010001010" => data <= "000000";
				when "001100100010001011" => data <= "000000";
				when "001100100010001100" => data <= "000000";
				when "001100100010001101" => data <= "000000";
				when "001100100010001110" => data <= "000000";
				when "001100100010001111" => data <= "000000";
				when "001100100010010000" => data <= "000000";
				when "001100100010010001" => data <= "000000";
				when "001100100010010010" => data <= "000000";
				when "001100100010010011" => data <= "000000";
				when "001100100010010100" => data <= "000000";
				when "001100100010010101" => data <= "000000";
				when "001100100010010110" => data <= "000000";
				when "001100100010010111" => data <= "000000";
				when "001100100010011000" => data <= "000000";
				when "001100100010011001" => data <= "000000";
				when "001100100010011010" => data <= "000000";
				when "001100100010011011" => data <= "000000";
				when "001100100010011100" => data <= "000000";
				when "001100100010011101" => data <= "000000";
				when "001100100010011110" => data <= "000000";
				when "001100100010011111" => data <= "000000";
				when "001100101000000000" => data <= "000000";
				when "001100101000000001" => data <= "000000";
				when "001100101000000010" => data <= "000000";
				when "001100101000000011" => data <= "000000";
				when "001100101000000100" => data <= "000000";
				when "001100101000000101" => data <= "000000";
				when "001100101000000110" => data <= "000000";
				when "001100101000000111" => data <= "000000";
				when "001100101000001000" => data <= "000000";
				when "001100101000001001" => data <= "000000";
				when "001100101000001010" => data <= "000000";
				when "001100101000001011" => data <= "000000";
				when "001100101000001100" => data <= "000000";
				when "001100101000001101" => data <= "000000";
				when "001100101000001110" => data <= "000000";
				when "001100101000001111" => data <= "000000";
				when "001100101000010000" => data <= "000000";
				when "001100101000010001" => data <= "000000";
				when "001100101000010010" => data <= "000000";
				when "001100101000010011" => data <= "000000";
				when "001100101000010100" => data <= "000000";
				when "001100101000010101" => data <= "000000";
				when "001100101000010110" => data <= "000000";
				when "001100101000010111" => data <= "000000";
				when "001100101000011000" => data <= "000000";
				when "001100101000011001" => data <= "000000";
				when "001100101000011010" => data <= "000000";
				when "001100101000011011" => data <= "000000";
				when "001100101000011100" => data <= "000000";
				when "001100101000011101" => data <= "000000";
				when "001100101000011110" => data <= "000000";
				when "001100101000011111" => data <= "000000";
				when "001100101000100000" => data <= "000000";
				when "001100101000100001" => data <= "000000";
				when "001100101000100010" => data <= "000000";
				when "001100101000100011" => data <= "000000";
				when "001100101000100100" => data <= "000000";
				when "001100101000100101" => data <= "000000";
				when "001100101000100110" => data <= "000000";
				when "001100101000100111" => data <= "000000";
				when "001100101000101000" => data <= "000000";
				when "001100101000101001" => data <= "000000";
				when "001100101000101010" => data <= "000000";
				when "001100101000101011" => data <= "000000";
				when "001100101000101100" => data <= "000000";
				when "001100101000101101" => data <= "000000";
				when "001100101000101110" => data <= "000000";
				when "001100101000101111" => data <= "000000";
				when "001100101000110000" => data <= "000000";
				when "001100101000110001" => data <= "000000";
				when "001100101000110010" => data <= "000000";
				when "001100101000110011" => data <= "000000";
				when "001100101000110100" => data <= "000000";
				when "001100101000110101" => data <= "000000";
				when "001100101000110110" => data <= "000000";
				when "001100101000110111" => data <= "000000";
				when "001100101000111000" => data <= "000000";
				when "001100101000111001" => data <= "000000";
				when "001100101000111010" => data <= "000000";
				when "001100101000111011" => data <= "000000";
				when "001100101000111100" => data <= "000000";
				when "001100101000111101" => data <= "000000";
				when "001100101000111110" => data <= "000000";
				when "001100101000111111" => data <= "000000";
				when "001100101001000000" => data <= "000000";
				when "001100101001000001" => data <= "000000";
				when "001100101001000010" => data <= "000000";
				when "001100101001000011" => data <= "000000";
				when "001100101001000100" => data <= "000000";
				when "001100101001000101" => data <= "000000";
				when "001100101001000110" => data <= "000000";
				when "001100101001000111" => data <= "000000";
				when "001100101001001000" => data <= "000000";
				when "001100101001001001" => data <= "000000";
				when "001100101001001010" => data <= "000000";
				when "001100101001001011" => data <= "000000";
				when "001100101001001100" => data <= "000000";
				when "001100101001001101" => data <= "000000";
				when "001100101001001110" => data <= "000000";
				when "001100101001001111" => data <= "000000";
				when "001100101001010000" => data <= "000000";
				when "001100101001010001" => data <= "000000";
				when "001100101001010010" => data <= "000000";
				when "001100101001010011" => data <= "000000";
				when "001100101001010100" => data <= "000000";
				when "001100101001010101" => data <= "000000";
				when "001100101001010110" => data <= "000000";
				when "001100101001010111" => data <= "000000";
				when "001100101001011000" => data <= "000000";
				when "001100101001011001" => data <= "000000";
				when "001100101001011010" => data <= "000000";
				when "001100101001011011" => data <= "000000";
				when "001100101001011100" => data <= "000000";
				when "001100101001011101" => data <= "000000";
				when "001100101001011110" => data <= "000000";
				when "001100101001011111" => data <= "000000";
				when "001100101001100000" => data <= "000000";
				when "001100101001100001" => data <= "000000";
				when "001100101001100010" => data <= "000000";
				when "001100101001100011" => data <= "000000";
				when "001100101001100100" => data <= "000000";
				when "001100101001100101" => data <= "000000";
				when "001100101001100110" => data <= "000000";
				when "001100101001100111" => data <= "000000";
				when "001100101001101000" => data <= "000000";
				when "001100101001101001" => data <= "000000";
				when "001100101001101010" => data <= "000000";
				when "001100101001101011" => data <= "000000";
				when "001100101001101100" => data <= "000000";
				when "001100101001101101" => data <= "000000";
				when "001100101001101110" => data <= "000000";
				when "001100101001101111" => data <= "000000";
				when "001100101001110000" => data <= "000000";
				when "001100101001110001" => data <= "000000";
				when "001100101001110010" => data <= "000000";
				when "001100101001110011" => data <= "000000";
				when "001100101001110100" => data <= "000000";
				when "001100101001110101" => data <= "000000";
				when "001100101001110110" => data <= "000000";
				when "001100101001110111" => data <= "000000";
				when "001100101001111000" => data <= "000000";
				when "001100101001111001" => data <= "000000";
				when "001100101001111010" => data <= "000000";
				when "001100101001111011" => data <= "000000";
				when "001100101001111100" => data <= "000000";
				when "001100101001111101" => data <= "000000";
				when "001100101001111110" => data <= "000000";
				when "001100101001111111" => data <= "000000";
				when "001100101010000000" => data <= "000000";
				when "001100101010000001" => data <= "000000";
				when "001100101010000010" => data <= "000000";
				when "001100101010000011" => data <= "000000";
				when "001100101010000100" => data <= "000000";
				when "001100101010000101" => data <= "000000";
				when "001100101010000110" => data <= "000000";
				when "001100101010000111" => data <= "000000";
				when "001100101010001000" => data <= "000000";
				when "001100101010001001" => data <= "000000";
				when "001100101010001010" => data <= "000000";
				when "001100101010001011" => data <= "000000";
				when "001100101010001100" => data <= "000000";
				when "001100101010001101" => data <= "000000";
				when "001100101010001110" => data <= "000000";
				when "001100101010001111" => data <= "000000";
				when "001100101010010000" => data <= "000000";
				when "001100101010010001" => data <= "000000";
				when "001100101010010010" => data <= "000000";
				when "001100101010010011" => data <= "000000";
				when "001100101010010100" => data <= "000000";
				when "001100101010010101" => data <= "000000";
				when "001100101010010110" => data <= "000000";
				when "001100101010010111" => data <= "000000";
				when "001100101010011000" => data <= "000000";
				when "001100101010011001" => data <= "000000";
				when "001100101010011010" => data <= "000000";
				when "001100101010011011" => data <= "000000";
				when "001100101010011100" => data <= "000000";
				when "001100101010011101" => data <= "000000";
				when "001100101010011110" => data <= "000000";
				when "001100101010011111" => data <= "000000";
				when "001100110000000000" => data <= "000000";
				when "001100110000000001" => data <= "000000";
				when "001100110000000010" => data <= "000000";
				when "001100110000000011" => data <= "000000";
				when "001100110000000100" => data <= "000000";
				when "001100110000000101" => data <= "000000";
				when "001100110000000110" => data <= "000000";
				when "001100110000000111" => data <= "000000";
				when "001100110000001000" => data <= "000000";
				when "001100110000001001" => data <= "000000";
				when "001100110000001010" => data <= "000000";
				when "001100110000001011" => data <= "000000";
				when "001100110000001100" => data <= "000000";
				when "001100110000001101" => data <= "000000";
				when "001100110000001110" => data <= "000000";
				when "001100110000001111" => data <= "000000";
				when "001100110000010000" => data <= "000000";
				when "001100110000010001" => data <= "000000";
				when "001100110000010010" => data <= "000000";
				when "001100110000010011" => data <= "000000";
				when "001100110000010100" => data <= "000000";
				when "001100110000010101" => data <= "000000";
				when "001100110000010110" => data <= "000000";
				when "001100110000010111" => data <= "000000";
				when "001100110000011000" => data <= "000000";
				when "001100110000011001" => data <= "000000";
				when "001100110000011010" => data <= "000000";
				when "001100110000011011" => data <= "000000";
				when "001100110000011100" => data <= "000000";
				when "001100110000011101" => data <= "000000";
				when "001100110000011110" => data <= "000000";
				when "001100110000011111" => data <= "000000";
				when "001100110000100000" => data <= "000000";
				when "001100110000100001" => data <= "000000";
				when "001100110000100010" => data <= "000000";
				when "001100110000100011" => data <= "000000";
				when "001100110000100100" => data <= "000000";
				when "001100110000100101" => data <= "000000";
				when "001100110000100110" => data <= "000000";
				when "001100110000100111" => data <= "000000";
				when "001100110000101000" => data <= "000000";
				when "001100110000101001" => data <= "000000";
				when "001100110000101010" => data <= "000000";
				when "001100110000101011" => data <= "000000";
				when "001100110000101100" => data <= "000000";
				when "001100110000101101" => data <= "000000";
				when "001100110000101110" => data <= "000000";
				when "001100110000101111" => data <= "000000";
				when "001100110000110000" => data <= "000000";
				when "001100110000110001" => data <= "000000";
				when "001100110000110010" => data <= "000000";
				when "001100110000110011" => data <= "000000";
				when "001100110000110100" => data <= "000000";
				when "001100110000110101" => data <= "000000";
				when "001100110000110110" => data <= "000000";
				when "001100110000110111" => data <= "000000";
				when "001100110000111000" => data <= "000000";
				when "001100110000111001" => data <= "000000";
				when "001100110000111010" => data <= "000000";
				when "001100110000111011" => data <= "000000";
				when "001100110000111100" => data <= "000000";
				when "001100110000111101" => data <= "000000";
				when "001100110000111110" => data <= "000000";
				when "001100110000111111" => data <= "000000";
				when "001100110001000000" => data <= "000000";
				when "001100110001000001" => data <= "000000";
				when "001100110001000010" => data <= "000000";
				when "001100110001000011" => data <= "000000";
				when "001100110001000100" => data <= "000000";
				when "001100110001000101" => data <= "000000";
				when "001100110001000110" => data <= "000000";
				when "001100110001000111" => data <= "000000";
				when "001100110001001000" => data <= "000000";
				when "001100110001001001" => data <= "000000";
				when "001100110001001010" => data <= "000000";
				when "001100110001001011" => data <= "000000";
				when "001100110001001100" => data <= "000000";
				when "001100110001001101" => data <= "000000";
				when "001100110001001110" => data <= "000000";
				when "001100110001001111" => data <= "000000";
				when "001100110001010000" => data <= "000000";
				when "001100110001010001" => data <= "000000";
				when "001100110001010010" => data <= "000000";
				when "001100110001010011" => data <= "000000";
				when "001100110001010100" => data <= "000000";
				when "001100110001010101" => data <= "000000";
				when "001100110001010110" => data <= "000000";
				when "001100110001010111" => data <= "000000";
				when "001100110001011000" => data <= "000000";
				when "001100110001011001" => data <= "000000";
				when "001100110001011010" => data <= "000000";
				when "001100110001011011" => data <= "000000";
				when "001100110001011100" => data <= "000000";
				when "001100110001011101" => data <= "000000";
				when "001100110001011110" => data <= "000000";
				when "001100110001011111" => data <= "000000";
				when "001100110001100000" => data <= "000000";
				when "001100110001100001" => data <= "000000";
				when "001100110001100010" => data <= "000000";
				when "001100110001100011" => data <= "000000";
				when "001100110001100100" => data <= "000000";
				when "001100110001100101" => data <= "000000";
				when "001100110001100110" => data <= "000000";
				when "001100110001100111" => data <= "000000";
				when "001100110001101000" => data <= "000000";
				when "001100110001101001" => data <= "000000";
				when "001100110001101010" => data <= "000000";
				when "001100110001101011" => data <= "000000";
				when "001100110001101100" => data <= "000000";
				when "001100110001101101" => data <= "000000";
				when "001100110001101110" => data <= "000000";
				when "001100110001101111" => data <= "000000";
				when "001100110001110000" => data <= "000000";
				when "001100110001110001" => data <= "000000";
				when "001100110001110010" => data <= "000000";
				when "001100110001110011" => data <= "000000";
				when "001100110001110100" => data <= "000000";
				when "001100110001110101" => data <= "000000";
				when "001100110001110110" => data <= "000000";
				when "001100110001110111" => data <= "000000";
				when "001100110001111000" => data <= "000000";
				when "001100110001111001" => data <= "000000";
				when "001100110001111010" => data <= "000000";
				when "001100110001111011" => data <= "000000";
				when "001100110001111100" => data <= "000000";
				when "001100110001111101" => data <= "000000";
				when "001100110001111110" => data <= "000000";
				when "001100110001111111" => data <= "000000";
				when "001100110010000000" => data <= "000000";
				when "001100110010000001" => data <= "000000";
				when "001100110010000010" => data <= "000000";
				when "001100110010000011" => data <= "000000";
				when "001100110010000100" => data <= "000000";
				when "001100110010000101" => data <= "000000";
				when "001100110010000110" => data <= "000000";
				when "001100110010000111" => data <= "000000";
				when "001100110010001000" => data <= "000000";
				when "001100110010001001" => data <= "000000";
				when "001100110010001010" => data <= "000000";
				when "001100110010001011" => data <= "000000";
				when "001100110010001100" => data <= "000000";
				when "001100110010001101" => data <= "000000";
				when "001100110010001110" => data <= "000000";
				when "001100110010001111" => data <= "000000";
				when "001100110010010000" => data <= "000000";
				when "001100110010010001" => data <= "000000";
				when "001100110010010010" => data <= "000000";
				when "001100110010010011" => data <= "000000";
				when "001100110010010100" => data <= "000000";
				when "001100110010010101" => data <= "000000";
				when "001100110010010110" => data <= "000000";
				when "001100110010010111" => data <= "000000";
				when "001100110010011000" => data <= "000000";
				when "001100110010011001" => data <= "000000";
				when "001100110010011010" => data <= "000000";
				when "001100110010011011" => data <= "000000";
				when "001100110010011100" => data <= "000000";
				when "001100110010011101" => data <= "000000";
				when "001100110010011110" => data <= "000000";
				when "001100110010011111" => data <= "000000";
				when "001100111000000000" => data <= "000000";
				when "001100111000000001" => data <= "000000";
				when "001100111000000010" => data <= "000000";
				when "001100111000000011" => data <= "000000";
				when "001100111000000100" => data <= "000000";
				when "001100111000000101" => data <= "000000";
				when "001100111000000110" => data <= "000000";
				when "001100111000000111" => data <= "000000";
				when "001100111000001000" => data <= "000000";
				when "001100111000001001" => data <= "000000";
				when "001100111000001010" => data <= "000000";
				when "001100111000001011" => data <= "000000";
				when "001100111000001100" => data <= "000000";
				when "001100111000001101" => data <= "000000";
				when "001100111000001110" => data <= "000000";
				when "001100111000001111" => data <= "000000";
				when "001100111000010000" => data <= "000000";
				when "001100111000010001" => data <= "000000";
				when "001100111000010010" => data <= "000000";
				when "001100111000010011" => data <= "000000";
				when "001100111000010100" => data <= "000000";
				when "001100111000010101" => data <= "000000";
				when "001100111000010110" => data <= "000000";
				when "001100111000010111" => data <= "000000";
				when "001100111000011000" => data <= "000000";
				when "001100111000011001" => data <= "000000";
				when "001100111000011010" => data <= "000000";
				when "001100111000011011" => data <= "000000";
				when "001100111000011100" => data <= "000000";
				when "001100111000011101" => data <= "000000";
				when "001100111000011110" => data <= "000000";
				when "001100111000011111" => data <= "000000";
				when "001100111000100000" => data <= "000000";
				when "001100111000100001" => data <= "000000";
				when "001100111000100010" => data <= "000000";
				when "001100111000100011" => data <= "000000";
				when "001100111000100100" => data <= "000000";
				when "001100111000100101" => data <= "000000";
				when "001100111000100110" => data <= "000000";
				when "001100111000100111" => data <= "000000";
				when "001100111000101000" => data <= "000000";
				when "001100111000101001" => data <= "000000";
				when "001100111000101010" => data <= "000000";
				when "001100111000101011" => data <= "000000";
				when "001100111000101100" => data <= "000000";
				when "001100111000101101" => data <= "000000";
				when "001100111000101110" => data <= "000000";
				when "001100111000101111" => data <= "000000";
				when "001100111000110000" => data <= "000000";
				when "001100111000110001" => data <= "000000";
				when "001100111000110010" => data <= "000000";
				when "001100111000110011" => data <= "000000";
				when "001100111000110100" => data <= "000000";
				when "001100111000110101" => data <= "000000";
				when "001100111000110110" => data <= "000000";
				when "001100111000110111" => data <= "000000";
				when "001100111000111000" => data <= "000000";
				when "001100111000111001" => data <= "000000";
				when "001100111000111010" => data <= "000000";
				when "001100111000111011" => data <= "000000";
				when "001100111000111100" => data <= "000000";
				when "001100111000111101" => data <= "000000";
				when "001100111000111110" => data <= "000000";
				when "001100111000111111" => data <= "000000";
				when "001100111001000000" => data <= "000000";
				when "001100111001000001" => data <= "000000";
				when "001100111001000010" => data <= "000000";
				when "001100111001000011" => data <= "000000";
				when "001100111001000100" => data <= "000000";
				when "001100111001000101" => data <= "000000";
				when "001100111001000110" => data <= "000000";
				when "001100111001000111" => data <= "000000";
				when "001100111001001000" => data <= "000000";
				when "001100111001001001" => data <= "000000";
				when "001100111001001010" => data <= "000000";
				when "001100111001001011" => data <= "000000";
				when "001100111001001100" => data <= "000000";
				when "001100111001001101" => data <= "000000";
				when "001100111001001110" => data <= "000000";
				when "001100111001001111" => data <= "000000";
				when "001100111001010000" => data <= "000000";
				when "001100111001010001" => data <= "000000";
				when "001100111001010010" => data <= "000000";
				when "001100111001010011" => data <= "000000";
				when "001100111001010100" => data <= "000000";
				when "001100111001010101" => data <= "000000";
				when "001100111001010110" => data <= "000000";
				when "001100111001010111" => data <= "000000";
				when "001100111001011000" => data <= "000000";
				when "001100111001011001" => data <= "000000";
				when "001100111001011010" => data <= "000000";
				when "001100111001011011" => data <= "000000";
				when "001100111001011100" => data <= "000000";
				when "001100111001011101" => data <= "000000";
				when "001100111001011110" => data <= "000000";
				when "001100111001011111" => data <= "000000";
				when "001100111001100000" => data <= "000000";
				when "001100111001100001" => data <= "000000";
				when "001100111001100010" => data <= "000000";
				when "001100111001100011" => data <= "000000";
				when "001100111001100100" => data <= "000000";
				when "001100111001100101" => data <= "000000";
				when "001100111001100110" => data <= "000000";
				when "001100111001100111" => data <= "000000";
				when "001100111001101000" => data <= "000000";
				when "001100111001101001" => data <= "000000";
				when "001100111001101010" => data <= "000000";
				when "001100111001101011" => data <= "000000";
				when "001100111001101100" => data <= "000000";
				when "001100111001101101" => data <= "000000";
				when "001100111001101110" => data <= "000000";
				when "001100111001101111" => data <= "000000";
				when "001100111001110000" => data <= "000000";
				when "001100111001110001" => data <= "000000";
				when "001100111001110010" => data <= "000000";
				when "001100111001110011" => data <= "000000";
				when "001100111001110100" => data <= "000000";
				when "001100111001110101" => data <= "000000";
				when "001100111001110110" => data <= "000000";
				when "001100111001110111" => data <= "000000";
				when "001100111001111000" => data <= "000000";
				when "001100111001111001" => data <= "000000";
				when "001100111001111010" => data <= "000000";
				when "001100111001111011" => data <= "000000";
				when "001100111001111100" => data <= "000000";
				when "001100111001111101" => data <= "000000";
				when "001100111001111110" => data <= "000000";
				when "001100111001111111" => data <= "000000";
				when "001100111010000000" => data <= "000000";
				when "001100111010000001" => data <= "000000";
				when "001100111010000010" => data <= "000000";
				when "001100111010000011" => data <= "000000";
				when "001100111010000100" => data <= "000000";
				when "001100111010000101" => data <= "000000";
				when "001100111010000110" => data <= "000000";
				when "001100111010000111" => data <= "000000";
				when "001100111010001000" => data <= "000000";
				when "001100111010001001" => data <= "000000";
				when "001100111010001010" => data <= "000000";
				when "001100111010001011" => data <= "000000";
				when "001100111010001100" => data <= "000000";
				when "001100111010001101" => data <= "000000";
				when "001100111010001110" => data <= "000000";
				when "001100111010001111" => data <= "000000";
				when "001100111010010000" => data <= "000000";
				when "001100111010010001" => data <= "000000";
				when "001100111010010010" => data <= "000000";
				when "001100111010010011" => data <= "000000";
				when "001100111010010100" => data <= "000000";
				when "001100111010010101" => data <= "000000";
				when "001100111010010110" => data <= "000000";
				when "001100111010010111" => data <= "000000";
				when "001100111010011000" => data <= "000000";
				when "001100111010011001" => data <= "000000";
				when "001100111010011010" => data <= "000000";
				when "001100111010011011" => data <= "000000";
				when "001100111010011100" => data <= "000000";
				when "001100111010011101" => data <= "000000";
				when "001100111010011110" => data <= "000000";
				when "001100111010011111" => data <= "000000";
				when "001101000000000000" => data <= "000000";
				when "001101000000000001" => data <= "000000";
				when "001101000000000010" => data <= "000000";
				when "001101000000000011" => data <= "000000";
				when "001101000000000100" => data <= "000000";
				when "001101000000000101" => data <= "000000";
				when "001101000000000110" => data <= "000000";
				when "001101000000000111" => data <= "000000";
				when "001101000000001000" => data <= "000000";
				when "001101000000001001" => data <= "000000";
				when "001101000000001010" => data <= "000000";
				when "001101000000001011" => data <= "000000";
				when "001101000000001100" => data <= "000000";
				when "001101000000001101" => data <= "000000";
				when "001101000000001110" => data <= "000000";
				when "001101000000001111" => data <= "000000";
				when "001101000000010000" => data <= "000000";
				when "001101000000010001" => data <= "000000";
				when "001101000000010010" => data <= "000000";
				when "001101000000010011" => data <= "000000";
				when "001101000000010100" => data <= "000000";
				when "001101000000010101" => data <= "000000";
				when "001101000000010110" => data <= "000000";
				when "001101000000010111" => data <= "000000";
				when "001101000000011000" => data <= "000000";
				when "001101000000011001" => data <= "000000";
				when "001101000000011010" => data <= "000000";
				when "001101000000011011" => data <= "000000";
				when "001101000000011100" => data <= "000000";
				when "001101000000011101" => data <= "000000";
				when "001101000000011110" => data <= "000000";
				when "001101000000011111" => data <= "000000";
				when "001101000000100000" => data <= "000000";
				when "001101000000100001" => data <= "000000";
				when "001101000000100010" => data <= "000000";
				when "001101000000100011" => data <= "000000";
				when "001101000000100100" => data <= "000000";
				when "001101000000100101" => data <= "000000";
				when "001101000000100110" => data <= "000000";
				when "001101000000100111" => data <= "000000";
				when "001101000000101000" => data <= "000000";
				when "001101000000101001" => data <= "000000";
				when "001101000000101010" => data <= "000000";
				when "001101000000101011" => data <= "000000";
				when "001101000000101100" => data <= "000000";
				when "001101000000101101" => data <= "000000";
				when "001101000000101110" => data <= "000000";
				when "001101000000101111" => data <= "000000";
				when "001101000000110000" => data <= "000000";
				when "001101000000110001" => data <= "000000";
				when "001101000000110010" => data <= "000000";
				when "001101000000110011" => data <= "000000";
				when "001101000000110100" => data <= "000000";
				when "001101000000110101" => data <= "000000";
				when "001101000000110110" => data <= "000000";
				when "001101000000110111" => data <= "000000";
				when "001101000000111000" => data <= "000000";
				when "001101000000111001" => data <= "000000";
				when "001101000000111010" => data <= "000000";
				when "001101000000111011" => data <= "000000";
				when "001101000000111100" => data <= "000000";
				when "001101000000111101" => data <= "000000";
				when "001101000000111110" => data <= "000000";
				when "001101000000111111" => data <= "000000";
				when "001101000001000000" => data <= "000000";
				when "001101000001000001" => data <= "000000";
				when "001101000001000010" => data <= "000000";
				when "001101000001000011" => data <= "000000";
				when "001101000001000100" => data <= "000000";
				when "001101000001000101" => data <= "000000";
				when "001101000001000110" => data <= "000000";
				when "001101000001000111" => data <= "000000";
				when "001101000001001000" => data <= "000000";
				when "001101000001001001" => data <= "000000";
				when "001101000001001010" => data <= "000000";
				when "001101000001001011" => data <= "000000";
				when "001101000001001100" => data <= "000000";
				when "001101000001001101" => data <= "000000";
				when "001101000001001110" => data <= "000000";
				when "001101000001001111" => data <= "000000";
				when "001101000001010000" => data <= "000000";
				when "001101000001010001" => data <= "000000";
				when "001101000001010010" => data <= "000000";
				when "001101000001010011" => data <= "000000";
				when "001101000001010100" => data <= "000000";
				when "001101000001010101" => data <= "000000";
				when "001101000001010110" => data <= "000000";
				when "001101000001010111" => data <= "000000";
				when "001101000001011000" => data <= "000000";
				when "001101000001011001" => data <= "000000";
				when "001101000001011010" => data <= "000000";
				when "001101000001011011" => data <= "000000";
				when "001101000001011100" => data <= "000000";
				when "001101000001011101" => data <= "000000";
				when "001101000001011110" => data <= "000000";
				when "001101000001011111" => data <= "000000";
				when "001101000001100000" => data <= "000000";
				when "001101000001100001" => data <= "000000";
				when "001101000001100010" => data <= "000000";
				when "001101000001100011" => data <= "000000";
				when "001101000001100100" => data <= "000000";
				when "001101000001100101" => data <= "000000";
				when "001101000001100110" => data <= "000000";
				when "001101000001100111" => data <= "000000";
				when "001101000001101000" => data <= "000000";
				when "001101000001101001" => data <= "000000";
				when "001101000001101010" => data <= "000000";
				when "001101000001101011" => data <= "000000";
				when "001101000001101100" => data <= "000000";
				when "001101000001101101" => data <= "000000";
				when "001101000001101110" => data <= "000000";
				when "001101000001101111" => data <= "000000";
				when "001101000001110000" => data <= "000000";
				when "001101000001110001" => data <= "000000";
				when "001101000001110010" => data <= "000000";
				when "001101000001110011" => data <= "000000";
				when "001101000001110100" => data <= "000000";
				when "001101000001110101" => data <= "000000";
				when "001101000001110110" => data <= "000000";
				when "001101000001110111" => data <= "000000";
				when "001101000001111000" => data <= "000000";
				when "001101000001111001" => data <= "000000";
				when "001101000001111010" => data <= "000000";
				when "001101000001111011" => data <= "000000";
				when "001101000001111100" => data <= "000000";
				when "001101000001111101" => data <= "000000";
				when "001101000001111110" => data <= "000000";
				when "001101000001111111" => data <= "000000";
				when "001101000010000000" => data <= "000000";
				when "001101000010000001" => data <= "000000";
				when "001101000010000010" => data <= "000000";
				when "001101000010000011" => data <= "000000";
				when "001101000010000100" => data <= "000000";
				when "001101000010000101" => data <= "000000";
				when "001101000010000110" => data <= "000000";
				when "001101000010000111" => data <= "000000";
				when "001101000010001000" => data <= "000000";
				when "001101000010001001" => data <= "000000";
				when "001101000010001010" => data <= "000000";
				when "001101000010001011" => data <= "000000";
				when "001101000010001100" => data <= "000000";
				when "001101000010001101" => data <= "000000";
				when "001101000010001110" => data <= "000000";
				when "001101000010001111" => data <= "000000";
				when "001101000010010000" => data <= "000000";
				when "001101000010010001" => data <= "000000";
				when "001101000010010010" => data <= "000000";
				when "001101000010010011" => data <= "000000";
				when "001101000010010100" => data <= "000000";
				when "001101000010010101" => data <= "000000";
				when "001101000010010110" => data <= "000000";
				when "001101000010010111" => data <= "000000";
				when "001101000010011000" => data <= "000000";
				when "001101000010011001" => data <= "000000";
				when "001101000010011010" => data <= "000000";
				when "001101000010011011" => data <= "000000";
				when "001101000010011100" => data <= "000000";
				when "001101000010011101" => data <= "000000";
				when "001101000010011110" => data <= "000000";
				when "001101000010011111" => data <= "000000";
				when "001101001000000000" => data <= "000000";
				when "001101001000000001" => data <= "000000";
				when "001101001000000010" => data <= "000000";
				when "001101001000000011" => data <= "000000";
				when "001101001000000100" => data <= "000000";
				when "001101001000000101" => data <= "000000";
				when "001101001000000110" => data <= "000000";
				when "001101001000000111" => data <= "000000";
				when "001101001000001000" => data <= "000000";
				when "001101001000001001" => data <= "000000";
				when "001101001000001010" => data <= "000000";
				when "001101001000001011" => data <= "000000";
				when "001101001000001100" => data <= "000000";
				when "001101001000001101" => data <= "000000";
				when "001101001000001110" => data <= "000000";
				when "001101001000001111" => data <= "000000";
				when "001101001000010000" => data <= "000000";
				when "001101001000010001" => data <= "000000";
				when "001101001000010010" => data <= "000000";
				when "001101001000010011" => data <= "000000";
				when "001101001000010100" => data <= "000000";
				when "001101001000010101" => data <= "000000";
				when "001101001000010110" => data <= "000000";
				when "001101001000010111" => data <= "000000";
				when "001101001000011000" => data <= "000000";
				when "001101001000011001" => data <= "000000";
				when "001101001000011010" => data <= "000000";
				when "001101001000011011" => data <= "000000";
				when "001101001000011100" => data <= "000000";
				when "001101001000011101" => data <= "000000";
				when "001101001000011110" => data <= "000000";
				when "001101001000011111" => data <= "000000";
				when "001101001000100000" => data <= "000000";
				when "001101001000100001" => data <= "000000";
				when "001101001000100010" => data <= "000000";
				when "001101001000100011" => data <= "000000";
				when "001101001000100100" => data <= "000000";
				when "001101001000100101" => data <= "000000";
				when "001101001000100110" => data <= "000000";
				when "001101001000100111" => data <= "000000";
				when "001101001000101000" => data <= "000000";
				when "001101001000101001" => data <= "000000";
				when "001101001000101010" => data <= "000000";
				when "001101001000101011" => data <= "000000";
				when "001101001000101100" => data <= "000000";
				when "001101001000101101" => data <= "000000";
				when "001101001000101110" => data <= "000000";
				when "001101001000101111" => data <= "000000";
				when "001101001000110000" => data <= "000000";
				when "001101001000110001" => data <= "000000";
				when "001101001000110010" => data <= "000000";
				when "001101001000110011" => data <= "000000";
				when "001101001000110100" => data <= "000000";
				when "001101001000110101" => data <= "000000";
				when "001101001000110110" => data <= "000000";
				when "001101001000110111" => data <= "000000";
				when "001101001000111000" => data <= "000000";
				when "001101001000111001" => data <= "000000";
				when "001101001000111010" => data <= "000000";
				when "001101001000111011" => data <= "000000";
				when "001101001000111100" => data <= "000000";
				when "001101001000111101" => data <= "000000";
				when "001101001000111110" => data <= "000000";
				when "001101001000111111" => data <= "000000";
				when "001101001001000000" => data <= "000000";
				when "001101001001000001" => data <= "000000";
				when "001101001001000010" => data <= "000000";
				when "001101001001000011" => data <= "000000";
				when "001101001001000100" => data <= "000000";
				when "001101001001000101" => data <= "000000";
				when "001101001001000110" => data <= "000000";
				when "001101001001000111" => data <= "000000";
				when "001101001001001000" => data <= "000000";
				when "001101001001001001" => data <= "000000";
				when "001101001001001010" => data <= "000000";
				when "001101001001001011" => data <= "000000";
				when "001101001001001100" => data <= "000000";
				when "001101001001001101" => data <= "000000";
				when "001101001001001110" => data <= "000000";
				when "001101001001001111" => data <= "000000";
				when "001101001001010000" => data <= "000000";
				when "001101001001010001" => data <= "000000";
				when "001101001001010010" => data <= "000000";
				when "001101001001010011" => data <= "000000";
				when "001101001001010100" => data <= "000000";
				when "001101001001010101" => data <= "000000";
				when "001101001001010110" => data <= "000000";
				when "001101001001010111" => data <= "000000";
				when "001101001001011000" => data <= "000000";
				when "001101001001011001" => data <= "000000";
				when "001101001001011010" => data <= "000000";
				when "001101001001011011" => data <= "000000";
				when "001101001001011100" => data <= "000000";
				when "001101001001011101" => data <= "000000";
				when "001101001001011110" => data <= "000000";
				when "001101001001011111" => data <= "000000";
				when "001101001001100000" => data <= "000000";
				when "001101001001100001" => data <= "000000";
				when "001101001001100010" => data <= "000000";
				when "001101001001100011" => data <= "000000";
				when "001101001001100100" => data <= "000000";
				when "001101001001100101" => data <= "000000";
				when "001101001001100110" => data <= "000000";
				when "001101001001100111" => data <= "000000";
				when "001101001001101000" => data <= "000000";
				when "001101001001101001" => data <= "000000";
				when "001101001001101010" => data <= "000000";
				when "001101001001101011" => data <= "000000";
				when "001101001001101100" => data <= "000000";
				when "001101001001101101" => data <= "000000";
				when "001101001001101110" => data <= "000000";
				when "001101001001101111" => data <= "000000";
				when "001101001001110000" => data <= "000000";
				when "001101001001110001" => data <= "000000";
				when "001101001001110010" => data <= "000000";
				when "001101001001110011" => data <= "000000";
				when "001101001001110100" => data <= "000000";
				when "001101001001110101" => data <= "000000";
				when "001101001001110110" => data <= "000000";
				when "001101001001110111" => data <= "000000";
				when "001101001001111000" => data <= "000000";
				when "001101001001111001" => data <= "000000";
				when "001101001001111010" => data <= "000000";
				when "001101001001111011" => data <= "000000";
				when "001101001001111100" => data <= "000000";
				when "001101001001111101" => data <= "000000";
				when "001101001001111110" => data <= "000000";
				when "001101001001111111" => data <= "000000";
				when "001101001010000000" => data <= "000000";
				when "001101001010000001" => data <= "000000";
				when "001101001010000010" => data <= "000000";
				when "001101001010000011" => data <= "000000";
				when "001101001010000100" => data <= "000000";
				when "001101001010000101" => data <= "000000";
				when "001101001010000110" => data <= "000000";
				when "001101001010000111" => data <= "000000";
				when "001101001010001000" => data <= "000000";
				when "001101001010001001" => data <= "000000";
				when "001101001010001010" => data <= "000000";
				when "001101001010001011" => data <= "000000";
				when "001101001010001100" => data <= "000000";
				when "001101001010001101" => data <= "000000";
				when "001101001010001110" => data <= "000000";
				when "001101001010001111" => data <= "000000";
				when "001101001010010000" => data <= "000000";
				when "001101001010010001" => data <= "000000";
				when "001101001010010010" => data <= "000000";
				when "001101001010010011" => data <= "000000";
				when "001101001010010100" => data <= "000000";
				when "001101001010010101" => data <= "000000";
				when "001101001010010110" => data <= "000000";
				when "001101001010010111" => data <= "000000";
				when "001101001010011000" => data <= "000000";
				when "001101001010011001" => data <= "000000";
				when "001101001010011010" => data <= "000000";
				when "001101001010011011" => data <= "000000";
				when "001101001010011100" => data <= "000000";
				when "001101001010011101" => data <= "000000";
				when "001101001010011110" => data <= "000000";
				when "001101001010011111" => data <= "000000";
				when "001101010000000000" => data <= "000000";
				when "001101010000000001" => data <= "000000";
				when "001101010000000010" => data <= "000000";
				when "001101010000000011" => data <= "000000";
				when "001101010000000100" => data <= "000000";
				when "001101010000000101" => data <= "000000";
				when "001101010000000110" => data <= "000000";
				when "001101010000000111" => data <= "000000";
				when "001101010000001000" => data <= "000000";
				when "001101010000001001" => data <= "000000";
				when "001101010000001010" => data <= "000000";
				when "001101010000001011" => data <= "000000";
				when "001101010000001100" => data <= "000000";
				when "001101010000001101" => data <= "000000";
				when "001101010000001110" => data <= "000000";
				when "001101010000001111" => data <= "000000";
				when "001101010000010000" => data <= "000000";
				when "001101010000010001" => data <= "000000";
				when "001101010000010010" => data <= "000000";
				when "001101010000010011" => data <= "000000";
				when "001101010000010100" => data <= "000000";
				when "001101010000010101" => data <= "000000";
				when "001101010000010110" => data <= "000000";
				when "001101010000010111" => data <= "000000";
				when "001101010000011000" => data <= "000000";
				when "001101010000011001" => data <= "000000";
				when "001101010000011010" => data <= "000000";
				when "001101010000011011" => data <= "000000";
				when "001101010000011100" => data <= "000000";
				when "001101010000011101" => data <= "000000";
				when "001101010000011110" => data <= "000000";
				when "001101010000011111" => data <= "000000";
				when "001101010000100000" => data <= "000000";
				when "001101010000100001" => data <= "000000";
				when "001101010000100010" => data <= "000000";
				when "001101010000100011" => data <= "000000";
				when "001101010000100100" => data <= "000000";
				when "001101010000100101" => data <= "000000";
				when "001101010000100110" => data <= "000000";
				when "001101010000100111" => data <= "000000";
				when "001101010000101000" => data <= "000000";
				when "001101010000101001" => data <= "000000";
				when "001101010000101010" => data <= "000000";
				when "001101010000101011" => data <= "000000";
				when "001101010000101100" => data <= "000000";
				when "001101010000101101" => data <= "000000";
				when "001101010000101110" => data <= "000000";
				when "001101010000101111" => data <= "000000";
				when "001101010000110000" => data <= "000000";
				when "001101010000110001" => data <= "000000";
				when "001101010000110010" => data <= "000000";
				when "001101010000110011" => data <= "000000";
				when "001101010000110100" => data <= "000000";
				when "001101010000110101" => data <= "000000";
				when "001101010000110110" => data <= "000000";
				when "001101010000110111" => data <= "000000";
				when "001101010000111000" => data <= "000000";
				when "001101010000111001" => data <= "000000";
				when "001101010000111010" => data <= "000000";
				when "001101010000111011" => data <= "000000";
				when "001101010000111100" => data <= "000000";
				when "001101010000111101" => data <= "000000";
				when "001101010000111110" => data <= "000000";
				when "001101010000111111" => data <= "000000";
				when "001101010001000000" => data <= "000000";
				when "001101010001000001" => data <= "000000";
				when "001101010001000010" => data <= "000000";
				when "001101010001000011" => data <= "000000";
				when "001101010001000100" => data <= "000000";
				when "001101010001000101" => data <= "000000";
				when "001101010001000110" => data <= "000000";
				when "001101010001000111" => data <= "000000";
				when "001101010001001000" => data <= "000000";
				when "001101010001001001" => data <= "000000";
				when "001101010001001010" => data <= "000000";
				when "001101010001001011" => data <= "000000";
				when "001101010001001100" => data <= "000000";
				when "001101010001001101" => data <= "000000";
				when "001101010001001110" => data <= "000000";
				when "001101010001001111" => data <= "000000";
				when "001101010001010000" => data <= "000000";
				when "001101010001010001" => data <= "000000";
				when "001101010001010010" => data <= "000000";
				when "001101010001010011" => data <= "000000";
				when "001101010001010100" => data <= "000000";
				when "001101010001010101" => data <= "000000";
				when "001101010001010110" => data <= "000000";
				when "001101010001010111" => data <= "000000";
				when "001101010001011000" => data <= "000000";
				when "001101010001011001" => data <= "000000";
				when "001101010001011010" => data <= "000000";
				when "001101010001011011" => data <= "000000";
				when "001101010001011100" => data <= "000000";
				when "001101010001011101" => data <= "000000";
				when "001101010001011110" => data <= "000000";
				when "001101010001011111" => data <= "000000";
				when "001101010001100000" => data <= "000000";
				when "001101010001100001" => data <= "000000";
				when "001101010001100010" => data <= "000000";
				when "001101010001100011" => data <= "000000";
				when "001101010001100100" => data <= "000000";
				when "001101010001100101" => data <= "000000";
				when "001101010001100110" => data <= "000000";
				when "001101010001100111" => data <= "000000";
				when "001101010001101000" => data <= "000000";
				when "001101010001101001" => data <= "000000";
				when "001101010001101010" => data <= "000000";
				when "001101010001101011" => data <= "000000";
				when "001101010001101100" => data <= "000000";
				when "001101010001101101" => data <= "000000";
				when "001101010001101110" => data <= "000000";
				when "001101010001101111" => data <= "000000";
				when "001101010001110000" => data <= "000000";
				when "001101010001110001" => data <= "000000";
				when "001101010001110010" => data <= "000000";
				when "001101010001110011" => data <= "000000";
				when "001101010001110100" => data <= "000000";
				when "001101010001110101" => data <= "000000";
				when "001101010001110110" => data <= "000000";
				when "001101010001110111" => data <= "000000";
				when "001101010001111000" => data <= "000000";
				when "001101010001111001" => data <= "000000";
				when "001101010001111010" => data <= "000000";
				when "001101010001111011" => data <= "000000";
				when "001101010001111100" => data <= "000000";
				when "001101010001111101" => data <= "000000";
				when "001101010001111110" => data <= "000000";
				when "001101010001111111" => data <= "000000";
				when "001101010010000000" => data <= "000000";
				when "001101010010000001" => data <= "000000";
				when "001101010010000010" => data <= "000000";
				when "001101010010000011" => data <= "000000";
				when "001101010010000100" => data <= "000000";
				when "001101010010000101" => data <= "000000";
				when "001101010010000110" => data <= "000000";
				when "001101010010000111" => data <= "000000";
				when "001101010010001000" => data <= "000000";
				when "001101010010001001" => data <= "000000";
				when "001101010010001010" => data <= "000000";
				when "001101010010001011" => data <= "000000";
				when "001101010010001100" => data <= "000000";
				when "001101010010001101" => data <= "000000";
				when "001101010010001110" => data <= "000000";
				when "001101010010001111" => data <= "000000";
				when "001101010010010000" => data <= "000000";
				when "001101010010010001" => data <= "000000";
				when "001101010010010010" => data <= "000000";
				when "001101010010010011" => data <= "000000";
				when "001101010010010100" => data <= "000000";
				when "001101010010010101" => data <= "000000";
				when "001101010010010110" => data <= "000000";
				when "001101010010010111" => data <= "000000";
				when "001101010010011000" => data <= "000000";
				when "001101010010011001" => data <= "000000";
				when "001101010010011010" => data <= "000000";
				when "001101010010011011" => data <= "000000";
				when "001101010010011100" => data <= "000000";
				when "001101010010011101" => data <= "000000";
				when "001101010010011110" => data <= "000000";
				when "001101010010011111" => data <= "000000";
				when "001101011000000000" => data <= "000000";
				when "001101011000000001" => data <= "000000";
				when "001101011000000010" => data <= "000000";
				when "001101011000000011" => data <= "000000";
				when "001101011000000100" => data <= "000000";
				when "001101011000000101" => data <= "000000";
				when "001101011000000110" => data <= "000000";
				when "001101011000000111" => data <= "000000";
				when "001101011000001000" => data <= "000000";
				when "001101011000001001" => data <= "000000";
				when "001101011000001010" => data <= "000000";
				when "001101011000001011" => data <= "000000";
				when "001101011000001100" => data <= "000000";
				when "001101011000001101" => data <= "000000";
				when "001101011000001110" => data <= "000000";
				when "001101011000001111" => data <= "000000";
				when "001101011000010000" => data <= "000000";
				when "001101011000010001" => data <= "000000";
				when "001101011000010010" => data <= "000000";
				when "001101011000010011" => data <= "000000";
				when "001101011000010100" => data <= "000000";
				when "001101011000010101" => data <= "000000";
				when "001101011000010110" => data <= "000000";
				when "001101011000010111" => data <= "000000";
				when "001101011000011000" => data <= "000000";
				when "001101011000011001" => data <= "000000";
				when "001101011000011010" => data <= "000000";
				when "001101011000011011" => data <= "000000";
				when "001101011000011100" => data <= "000000";
				when "001101011000011101" => data <= "000000";
				when "001101011000011110" => data <= "000000";
				when "001101011000011111" => data <= "000000";
				when "001101011000100000" => data <= "000000";
				when "001101011000100001" => data <= "000000";
				when "001101011000100010" => data <= "000000";
				when "001101011000100011" => data <= "000000";
				when "001101011000100100" => data <= "000000";
				when "001101011000100101" => data <= "000000";
				when "001101011000100110" => data <= "000000";
				when "001101011000100111" => data <= "000000";
				when "001101011000101000" => data <= "000000";
				when "001101011000101001" => data <= "000000";
				when "001101011000101010" => data <= "000000";
				when "001101011000101011" => data <= "000000";
				when "001101011000101100" => data <= "000000";
				when "001101011000101101" => data <= "000000";
				when "001101011000101110" => data <= "000000";
				when "001101011000101111" => data <= "000000";
				when "001101011000110000" => data <= "000000";
				when "001101011000110001" => data <= "000000";
				when "001101011000110010" => data <= "000000";
				when "001101011000110011" => data <= "000000";
				when "001101011000110100" => data <= "000000";
				when "001101011000110101" => data <= "000000";
				when "001101011000110110" => data <= "000000";
				when "001101011000110111" => data <= "000000";
				when "001101011000111000" => data <= "000000";
				when "001101011000111001" => data <= "000000";
				when "001101011000111010" => data <= "000000";
				when "001101011000111011" => data <= "000000";
				when "001101011000111100" => data <= "000000";
				when "001101011000111101" => data <= "000000";
				when "001101011000111110" => data <= "000000";
				when "001101011000111111" => data <= "000000";
				when "001101011001000000" => data <= "000000";
				when "001101011001000001" => data <= "000000";
				when "001101011001000010" => data <= "000000";
				when "001101011001000011" => data <= "000000";
				when "001101011001000100" => data <= "000000";
				when "001101011001000101" => data <= "000000";
				when "001101011001000110" => data <= "000000";
				when "001101011001000111" => data <= "000000";
				when "001101011001001000" => data <= "000000";
				when "001101011001001001" => data <= "000000";
				when "001101011001001010" => data <= "000000";
				when "001101011001001011" => data <= "000000";
				when "001101011001001100" => data <= "000000";
				when "001101011001001101" => data <= "000000";
				when "001101011001001110" => data <= "000000";
				when "001101011001001111" => data <= "000000";
				when "001101011001010000" => data <= "000000";
				when "001101011001010001" => data <= "000000";
				when "001101011001010010" => data <= "000000";
				when "001101011001010011" => data <= "000000";
				when "001101011001010100" => data <= "000000";
				when "001101011001010101" => data <= "000000";
				when "001101011001010110" => data <= "000000";
				when "001101011001010111" => data <= "000000";
				when "001101011001011000" => data <= "000000";
				when "001101011001011001" => data <= "000000";
				when "001101011001011010" => data <= "000000";
				when "001101011001011011" => data <= "000000";
				when "001101011001011100" => data <= "000000";
				when "001101011001011101" => data <= "000000";
				when "001101011001011110" => data <= "000000";
				when "001101011001011111" => data <= "000000";
				when "001101011001100000" => data <= "000000";
				when "001101011001100001" => data <= "000000";
				when "001101011001100010" => data <= "000000";
				when "001101011001100011" => data <= "000000";
				when "001101011001100100" => data <= "000000";
				when "001101011001100101" => data <= "000000";
				when "001101011001100110" => data <= "000000";
				when "001101011001100111" => data <= "000000";
				when "001101011001101000" => data <= "000000";
				when "001101011001101001" => data <= "000000";
				when "001101011001101010" => data <= "000000";
				when "001101011001101011" => data <= "000000";
				when "001101011001101100" => data <= "000000";
				when "001101011001101101" => data <= "000000";
				when "001101011001101110" => data <= "000000";
				when "001101011001101111" => data <= "000000";
				when "001101011001110000" => data <= "000000";
				when "001101011001110001" => data <= "000000";
				when "001101011001110010" => data <= "000000";
				when "001101011001110011" => data <= "000000";
				when "001101011001110100" => data <= "000000";
				when "001101011001110101" => data <= "000000";
				when "001101011001110110" => data <= "000000";
				when "001101011001110111" => data <= "000000";
				when "001101011001111000" => data <= "000000";
				when "001101011001111001" => data <= "000000";
				when "001101011001111010" => data <= "000000";
				when "001101011001111011" => data <= "000000";
				when "001101011001111100" => data <= "000000";
				when "001101011001111101" => data <= "000000";
				when "001101011001111110" => data <= "000000";
				when "001101011001111111" => data <= "000000";
				when "001101011010000000" => data <= "000000";
				when "001101011010000001" => data <= "000000";
				when "001101011010000010" => data <= "000000";
				when "001101011010000011" => data <= "000000";
				when "001101011010000100" => data <= "000000";
				when "001101011010000101" => data <= "000000";
				when "001101011010000110" => data <= "000000";
				when "001101011010000111" => data <= "000000";
				when "001101011010001000" => data <= "000000";
				when "001101011010001001" => data <= "000000";
				when "001101011010001010" => data <= "000000";
				when "001101011010001011" => data <= "000000";
				when "001101011010001100" => data <= "000000";
				when "001101011010001101" => data <= "000000";
				when "001101011010001110" => data <= "000000";
				when "001101011010001111" => data <= "000000";
				when "001101011010010000" => data <= "000000";
				when "001101011010010001" => data <= "000000";
				when "001101011010010010" => data <= "000000";
				when "001101011010010011" => data <= "000000";
				when "001101011010010100" => data <= "000000";
				when "001101011010010101" => data <= "000000";
				when "001101011010010110" => data <= "000000";
				when "001101011010010111" => data <= "000000";
				when "001101011010011000" => data <= "000000";
				when "001101011010011001" => data <= "000000";
				when "001101011010011010" => data <= "000000";
				when "001101011010011011" => data <= "000000";
				when "001101011010011100" => data <= "000000";
				when "001101011010011101" => data <= "000000";
				when "001101011010011110" => data <= "000000";
				when "001101011010011111" => data <= "000000";
				when "001101100000000000" => data <= "000000";
				when "001101100000000001" => data <= "000000";
				when "001101100000000010" => data <= "000000";
				when "001101100000000011" => data <= "000000";
				when "001101100000000100" => data <= "000000";
				when "001101100000000101" => data <= "000000";
				when "001101100000000110" => data <= "000000";
				when "001101100000000111" => data <= "000000";
				when "001101100000001000" => data <= "000000";
				when "001101100000001001" => data <= "000000";
				when "001101100000001010" => data <= "000000";
				when "001101100000001011" => data <= "000000";
				when "001101100000001100" => data <= "000000";
				when "001101100000001101" => data <= "000000";
				when "001101100000001110" => data <= "000000";
				when "001101100000001111" => data <= "000000";
				when "001101100000010000" => data <= "000000";
				when "001101100000010001" => data <= "000000";
				when "001101100000010010" => data <= "000000";
				when "001101100000010011" => data <= "000000";
				when "001101100000010100" => data <= "000000";
				when "001101100000010101" => data <= "000000";
				when "001101100000010110" => data <= "000000";
				when "001101100000010111" => data <= "000000";
				when "001101100000011000" => data <= "000000";
				when "001101100000011001" => data <= "000000";
				when "001101100000011010" => data <= "000000";
				when "001101100000011011" => data <= "000000";
				when "001101100000011100" => data <= "000000";
				when "001101100000011101" => data <= "000000";
				when "001101100000011110" => data <= "000000";
				when "001101100000011111" => data <= "000000";
				when "001101100000100000" => data <= "000000";
				when "001101100000100001" => data <= "000000";
				when "001101100000100010" => data <= "000000";
				when "001101100000100011" => data <= "000000";
				when "001101100000100100" => data <= "000000";
				when "001101100000100101" => data <= "000000";
				when "001101100000100110" => data <= "000000";
				when "001101100000100111" => data <= "000000";
				when "001101100000101000" => data <= "000000";
				when "001101100000101001" => data <= "000000";
				when "001101100000101010" => data <= "000000";
				when "001101100000101011" => data <= "000000";
				when "001101100000101100" => data <= "000000";
				when "001101100000101101" => data <= "000000";
				when "001101100000101110" => data <= "000000";
				when "001101100000101111" => data <= "000000";
				when "001101100000110000" => data <= "000000";
				when "001101100000110001" => data <= "000000";
				when "001101100000110010" => data <= "000000";
				when "001101100000110011" => data <= "000000";
				when "001101100000110100" => data <= "000000";
				when "001101100000110101" => data <= "000000";
				when "001101100000110110" => data <= "000000";
				when "001101100000110111" => data <= "000000";
				when "001101100000111000" => data <= "000000";
				when "001101100000111001" => data <= "000000";
				when "001101100000111010" => data <= "000000";
				when "001101100000111011" => data <= "000000";
				when "001101100000111100" => data <= "000000";
				when "001101100000111101" => data <= "000000";
				when "001101100000111110" => data <= "000000";
				when "001101100000111111" => data <= "000000";
				when "001101100001000000" => data <= "000000";
				when "001101100001000001" => data <= "000000";
				when "001101100001000010" => data <= "000000";
				when "001101100001000011" => data <= "000000";
				when "001101100001000100" => data <= "000000";
				when "001101100001000101" => data <= "000000";
				when "001101100001000110" => data <= "000000";
				when "001101100001000111" => data <= "000000";
				when "001101100001001000" => data <= "000000";
				when "001101100001001001" => data <= "000000";
				when "001101100001001010" => data <= "000000";
				when "001101100001001011" => data <= "000000";
				when "001101100001001100" => data <= "000000";
				when "001101100001001101" => data <= "000000";
				when "001101100001001110" => data <= "000000";
				when "001101100001001111" => data <= "000000";
				when "001101100001010000" => data <= "000000";
				when "001101100001010001" => data <= "000000";
				when "001101100001010010" => data <= "000000";
				when "001101100001010011" => data <= "000000";
				when "001101100001010100" => data <= "000000";
				when "001101100001010101" => data <= "000000";
				when "001101100001010110" => data <= "000000";
				when "001101100001010111" => data <= "000000";
				when "001101100001011000" => data <= "000000";
				when "001101100001011001" => data <= "000000";
				when "001101100001011010" => data <= "000000";
				when "001101100001011011" => data <= "000000";
				when "001101100001011100" => data <= "000000";
				when "001101100001011101" => data <= "000000";
				when "001101100001011110" => data <= "000000";
				when "001101100001011111" => data <= "000000";
				when "001101100001100000" => data <= "000000";
				when "001101100001100001" => data <= "000000";
				when "001101100001100010" => data <= "000000";
				when "001101100001100011" => data <= "000000";
				when "001101100001100100" => data <= "000000";
				when "001101100001100101" => data <= "000000";
				when "001101100001100110" => data <= "000000";
				when "001101100001100111" => data <= "000000";
				when "001101100001101000" => data <= "000000";
				when "001101100001101001" => data <= "000000";
				when "001101100001101010" => data <= "000000";
				when "001101100001101011" => data <= "000000";
				when "001101100001101100" => data <= "000000";
				when "001101100001101101" => data <= "000000";
				when "001101100001101110" => data <= "000000";
				when "001101100001101111" => data <= "000000";
				when "001101100001110000" => data <= "000000";
				when "001101100001110001" => data <= "000000";
				when "001101100001110010" => data <= "000000";
				when "001101100001110011" => data <= "000000";
				when "001101100001110100" => data <= "000000";
				when "001101100001110101" => data <= "000000";
				when "001101100001110110" => data <= "000000";
				when "001101100001110111" => data <= "000000";
				when "001101100001111000" => data <= "000000";
				when "001101100001111001" => data <= "000000";
				when "001101100001111010" => data <= "000000";
				when "001101100001111011" => data <= "000000";
				when "001101100001111100" => data <= "000000";
				when "001101100001111101" => data <= "000000";
				when "001101100001111110" => data <= "000000";
				when "001101100001111111" => data <= "000000";
				when "001101100010000000" => data <= "000000";
				when "001101100010000001" => data <= "000000";
				when "001101100010000010" => data <= "000000";
				when "001101100010000011" => data <= "000000";
				when "001101100010000100" => data <= "000000";
				when "001101100010000101" => data <= "000000";
				when "001101100010000110" => data <= "000000";
				when "001101100010000111" => data <= "000000";
				when "001101100010001000" => data <= "000000";
				when "001101100010001001" => data <= "000000";
				when "001101100010001010" => data <= "000000";
				when "001101100010001011" => data <= "000000";
				when "001101100010001100" => data <= "000000";
				when "001101100010001101" => data <= "000000";
				when "001101100010001110" => data <= "000000";
				when "001101100010001111" => data <= "000000";
				when "001101100010010000" => data <= "000000";
				when "001101100010010001" => data <= "000000";
				when "001101100010010010" => data <= "000000";
				when "001101100010010011" => data <= "000000";
				when "001101100010010100" => data <= "000000";
				when "001101100010010101" => data <= "000000";
				when "001101100010010110" => data <= "000000";
				when "001101100010010111" => data <= "000000";
				when "001101100010011000" => data <= "000000";
				when "001101100010011001" => data <= "000000";
				when "001101100010011010" => data <= "000000";
				when "001101100010011011" => data <= "000000";
				when "001101100010011100" => data <= "000000";
				when "001101100010011101" => data <= "000000";
				when "001101100010011110" => data <= "000000";
				when "001101100010011111" => data <= "000000";
				when "001101101000000000" => data <= "000000";
				when "001101101000000001" => data <= "000000";
				when "001101101000000010" => data <= "000000";
				when "001101101000000011" => data <= "000000";
				when "001101101000000100" => data <= "000000";
				when "001101101000000101" => data <= "000000";
				when "001101101000000110" => data <= "000000";
				when "001101101000000111" => data <= "000000";
				when "001101101000001000" => data <= "000000";
				when "001101101000001001" => data <= "000000";
				when "001101101000001010" => data <= "000000";
				when "001101101000001011" => data <= "000000";
				when "001101101000001100" => data <= "000000";
				when "001101101000001101" => data <= "000000";
				when "001101101000001110" => data <= "000000";
				when "001101101000001111" => data <= "000000";
				when "001101101000010000" => data <= "000000";
				when "001101101000010001" => data <= "000000";
				when "001101101000010010" => data <= "000000";
				when "001101101000010011" => data <= "000000";
				when "001101101000010100" => data <= "000000";
				when "001101101000010101" => data <= "000000";
				when "001101101000010110" => data <= "000000";
				when "001101101000010111" => data <= "000000";
				when "001101101000011000" => data <= "000000";
				when "001101101000011001" => data <= "000000";
				when "001101101000011010" => data <= "000000";
				when "001101101000011011" => data <= "000000";
				when "001101101000011100" => data <= "000000";
				when "001101101000011101" => data <= "000000";
				when "001101101000011110" => data <= "000000";
				when "001101101000011111" => data <= "000000";
				when "001101101000100000" => data <= "000000";
				when "001101101000100001" => data <= "000000";
				when "001101101000100010" => data <= "000000";
				when "001101101000100011" => data <= "000000";
				when "001101101000100100" => data <= "000000";
				when "001101101000100101" => data <= "000000";
				when "001101101000100110" => data <= "000000";
				when "001101101000100111" => data <= "000000";
				when "001101101000101000" => data <= "000000";
				when "001101101000101001" => data <= "000000";
				when "001101101000101010" => data <= "000000";
				when "001101101000101011" => data <= "000000";
				when "001101101000101100" => data <= "000000";
				when "001101101000101101" => data <= "000000";
				when "001101101000101110" => data <= "000000";
				when "001101101000101111" => data <= "000000";
				when "001101101000110000" => data <= "000000";
				when "001101101000110001" => data <= "000000";
				when "001101101000110010" => data <= "000000";
				when "001101101000110011" => data <= "000000";
				when "001101101000110100" => data <= "000000";
				when "001101101000110101" => data <= "000000";
				when "001101101000110110" => data <= "000000";
				when "001101101000110111" => data <= "000000";
				when "001101101000111000" => data <= "000000";
				when "001101101000111001" => data <= "000000";
				when "001101101000111010" => data <= "000000";
				when "001101101000111011" => data <= "000000";
				when "001101101000111100" => data <= "000000";
				when "001101101000111101" => data <= "000000";
				when "001101101000111110" => data <= "000000";
				when "001101101000111111" => data <= "000000";
				when "001101101001000000" => data <= "000000";
				when "001101101001000001" => data <= "000000";
				when "001101101001000010" => data <= "000000";
				when "001101101001000011" => data <= "000000";
				when "001101101001000100" => data <= "000000";
				when "001101101001000101" => data <= "000000";
				when "001101101001000110" => data <= "000000";
				when "001101101001000111" => data <= "000000";
				when "001101101001001000" => data <= "000000";
				when "001101101001001001" => data <= "000000";
				when "001101101001001010" => data <= "000000";
				when "001101101001001011" => data <= "000000";
				when "001101101001001100" => data <= "000000";
				when "001101101001001101" => data <= "000000";
				when "001101101001001110" => data <= "000000";
				when "001101101001001111" => data <= "000000";
				when "001101101001010000" => data <= "000000";
				when "001101101001010001" => data <= "000000";
				when "001101101001010010" => data <= "000000";
				when "001101101001010011" => data <= "000000";
				when "001101101001010100" => data <= "000000";
				when "001101101001010101" => data <= "000000";
				when "001101101001010110" => data <= "000000";
				when "001101101001010111" => data <= "000000";
				when "001101101001011000" => data <= "000000";
				when "001101101001011001" => data <= "000000";
				when "001101101001011010" => data <= "000000";
				when "001101101001011011" => data <= "000000";
				when "001101101001011100" => data <= "000000";
				when "001101101001011101" => data <= "000000";
				when "001101101001011110" => data <= "000000";
				when "001101101001011111" => data <= "000000";
				when "001101101001100000" => data <= "000000";
				when "001101101001100001" => data <= "000000";
				when "001101101001100010" => data <= "000000";
				when "001101101001100011" => data <= "000000";
				when "001101101001100100" => data <= "000000";
				when "001101101001100101" => data <= "000000";
				when "001101101001100110" => data <= "000000";
				when "001101101001100111" => data <= "000000";
				when "001101101001101000" => data <= "000000";
				when "001101101001101001" => data <= "000000";
				when "001101101001101010" => data <= "000000";
				when "001101101001101011" => data <= "000000";
				when "001101101001101100" => data <= "000000";
				when "001101101001101101" => data <= "000000";
				when "001101101001101110" => data <= "000000";
				when "001101101001101111" => data <= "000000";
				when "001101101001110000" => data <= "000000";
				when "001101101001110001" => data <= "000000";
				when "001101101001110010" => data <= "000000";
				when "001101101001110011" => data <= "000000";
				when "001101101001110100" => data <= "000000";
				when "001101101001110101" => data <= "000000";
				when "001101101001110110" => data <= "000000";
				when "001101101001110111" => data <= "000000";
				when "001101101001111000" => data <= "000000";
				when "001101101001111001" => data <= "000000";
				when "001101101001111010" => data <= "000000";
				when "001101101001111011" => data <= "000000";
				when "001101101001111100" => data <= "000000";
				when "001101101001111101" => data <= "000000";
				when "001101101001111110" => data <= "000000";
				when "001101101001111111" => data <= "000000";
				when "001101101010000000" => data <= "000000";
				when "001101101010000001" => data <= "000000";
				when "001101101010000010" => data <= "000000";
				when "001101101010000011" => data <= "000000";
				when "001101101010000100" => data <= "000000";
				when "001101101010000101" => data <= "000000";
				when "001101101010000110" => data <= "000000";
				when "001101101010000111" => data <= "000000";
				when "001101101010001000" => data <= "000000";
				when "001101101010001001" => data <= "000000";
				when "001101101010001010" => data <= "000000";
				when "001101101010001011" => data <= "000000";
				when "001101101010001100" => data <= "000000";
				when "001101101010001101" => data <= "000000";
				when "001101101010001110" => data <= "000000";
				when "001101101010001111" => data <= "000000";
				when "001101101010010000" => data <= "000000";
				when "001101101010010001" => data <= "000000";
				when "001101101010010010" => data <= "000000";
				when "001101101010010011" => data <= "000000";
				when "001101101010010100" => data <= "000000";
				when "001101101010010101" => data <= "000000";
				when "001101101010010110" => data <= "000000";
				when "001101101010010111" => data <= "000000";
				when "001101101010011000" => data <= "000000";
				when "001101101010011001" => data <= "000000";
				when "001101101010011010" => data <= "000000";
				when "001101101010011011" => data <= "000000";
				when "001101101010011100" => data <= "000000";
				when "001101101010011101" => data <= "000000";
				when "001101101010011110" => data <= "000000";
				when "001101101010011111" => data <= "000000";
				when "001101110000000000" => data <= "000000";
				when "001101110000000001" => data <= "000000";
				when "001101110000000010" => data <= "000000";
				when "001101110000000011" => data <= "000000";
				when "001101110000000100" => data <= "000000";
				when "001101110000000101" => data <= "000000";
				when "001101110000000110" => data <= "000000";
				when "001101110000000111" => data <= "000000";
				when "001101110000001000" => data <= "000000";
				when "001101110000001001" => data <= "000000";
				when "001101110000001010" => data <= "000000";
				when "001101110000001011" => data <= "000000";
				when "001101110000001100" => data <= "000000";
				when "001101110000001101" => data <= "000000";
				when "001101110000001110" => data <= "000000";
				when "001101110000001111" => data <= "000000";
				when "001101110000010000" => data <= "000000";
				when "001101110000010001" => data <= "000000";
				when "001101110000010010" => data <= "000000";
				when "001101110000010011" => data <= "000000";
				when "001101110000010100" => data <= "000000";
				when "001101110000010101" => data <= "000000";
				when "001101110000010110" => data <= "000000";
				when "001101110000010111" => data <= "000000";
				when "001101110000011000" => data <= "000000";
				when "001101110000011001" => data <= "000000";
				when "001101110000011010" => data <= "000000";
				when "001101110000011011" => data <= "000000";
				when "001101110000011100" => data <= "000000";
				when "001101110000011101" => data <= "000000";
				when "001101110000011110" => data <= "000000";
				when "001101110000011111" => data <= "000000";
				when "001101110000100000" => data <= "000000";
				when "001101110000100001" => data <= "000000";
				when "001101110000100010" => data <= "000000";
				when "001101110000100011" => data <= "000000";
				when "001101110000100100" => data <= "000000";
				when "001101110000100101" => data <= "000000";
				when "001101110000100110" => data <= "000000";
				when "001101110000100111" => data <= "000000";
				when "001101110000101000" => data <= "000000";
				when "001101110000101001" => data <= "000000";
				when "001101110000101010" => data <= "000000";
				when "001101110000101011" => data <= "000000";
				when "001101110000101100" => data <= "000000";
				when "001101110000101101" => data <= "000000";
				when "001101110000101110" => data <= "000000";
				when "001101110000101111" => data <= "000000";
				when "001101110000110000" => data <= "000000";
				when "001101110000110001" => data <= "000000";
				when "001101110000110010" => data <= "000000";
				when "001101110000110011" => data <= "000000";
				when "001101110000110100" => data <= "000000";
				when "001101110000110101" => data <= "000000";
				when "001101110000110110" => data <= "000000";
				when "001101110000110111" => data <= "000000";
				when "001101110000111000" => data <= "000000";
				when "001101110000111001" => data <= "000000";
				when "001101110000111010" => data <= "000000";
				when "001101110000111011" => data <= "000000";
				when "001101110000111100" => data <= "000000";
				when "001101110000111101" => data <= "000000";
				when "001101110000111110" => data <= "000000";
				when "001101110000111111" => data <= "000000";
				when "001101110001000000" => data <= "000000";
				when "001101110001000001" => data <= "000000";
				when "001101110001000010" => data <= "000000";
				when "001101110001000011" => data <= "000000";
				when "001101110001000100" => data <= "000000";
				when "001101110001000101" => data <= "000000";
				when "001101110001000110" => data <= "000000";
				when "001101110001000111" => data <= "000000";
				when "001101110001001000" => data <= "000000";
				when "001101110001001001" => data <= "000000";
				when "001101110001001010" => data <= "000000";
				when "001101110001001011" => data <= "000000";
				when "001101110001001100" => data <= "000000";
				when "001101110001001101" => data <= "000000";
				when "001101110001001110" => data <= "000000";
				when "001101110001001111" => data <= "000000";
				when "001101110001010000" => data <= "000000";
				when "001101110001010001" => data <= "000000";
				when "001101110001010010" => data <= "000000";
				when "001101110001010011" => data <= "000000";
				when "001101110001010100" => data <= "000000";
				when "001101110001010101" => data <= "000000";
				when "001101110001010110" => data <= "000000";
				when "001101110001010111" => data <= "000000";
				when "001101110001011000" => data <= "000000";
				when "001101110001011001" => data <= "000000";
				when "001101110001011010" => data <= "000000";
				when "001101110001011011" => data <= "000000";
				when "001101110001011100" => data <= "000000";
				when "001101110001011101" => data <= "000000";
				when "001101110001011110" => data <= "000000";
				when "001101110001011111" => data <= "000000";
				when "001101110001100000" => data <= "000000";
				when "001101110001100001" => data <= "000000";
				when "001101110001100010" => data <= "000000";
				when "001101110001100011" => data <= "000000";
				when "001101110001100100" => data <= "000000";
				when "001101110001100101" => data <= "000000";
				when "001101110001100110" => data <= "000000";
				when "001101110001100111" => data <= "000000";
				when "001101110001101000" => data <= "000000";
				when "001101110001101001" => data <= "000000";
				when "001101110001101010" => data <= "000000";
				when "001101110001101011" => data <= "000000";
				when "001101110001101100" => data <= "000000";
				when "001101110001101101" => data <= "000000";
				when "001101110001101110" => data <= "000000";
				when "001101110001101111" => data <= "000000";
				when "001101110001110000" => data <= "000000";
				when "001101110001110001" => data <= "000000";
				when "001101110001110010" => data <= "000000";
				when "001101110001110011" => data <= "000000";
				when "001101110001110100" => data <= "000000";
				when "001101110001110101" => data <= "000000";
				when "001101110001110110" => data <= "000000";
				when "001101110001110111" => data <= "000000";
				when "001101110001111000" => data <= "000000";
				when "001101110001111001" => data <= "000000";
				when "001101110001111010" => data <= "000000";
				when "001101110001111011" => data <= "000000";
				when "001101110001111100" => data <= "000000";
				when "001101110001111101" => data <= "000000";
				when "001101110001111110" => data <= "000000";
				when "001101110001111111" => data <= "000000";
				when "001101110010000000" => data <= "000000";
				when "001101110010000001" => data <= "000000";
				when "001101110010000010" => data <= "000000";
				when "001101110010000011" => data <= "000000";
				when "001101110010000100" => data <= "000000";
				when "001101110010000101" => data <= "000000";
				when "001101110010000110" => data <= "000000";
				when "001101110010000111" => data <= "000000";
				when "001101110010001000" => data <= "000000";
				when "001101110010001001" => data <= "000000";
				when "001101110010001010" => data <= "000000";
				when "001101110010001011" => data <= "000000";
				when "001101110010001100" => data <= "000000";
				when "001101110010001101" => data <= "000000";
				when "001101110010001110" => data <= "000000";
				when "001101110010001111" => data <= "000000";
				when "001101110010010000" => data <= "000000";
				when "001101110010010001" => data <= "000000";
				when "001101110010010010" => data <= "000000";
				when "001101110010010011" => data <= "000000";
				when "001101110010010100" => data <= "000000";
				when "001101110010010101" => data <= "000000";
				when "001101110010010110" => data <= "000000";
				when "001101110010010111" => data <= "000000";
				when "001101110010011000" => data <= "000000";
				when "001101110010011001" => data <= "000000";
				when "001101110010011010" => data <= "000000";
				when "001101110010011011" => data <= "000000";
				when "001101110010011100" => data <= "000000";
				when "001101110010011101" => data <= "000000";
				when "001101110010011110" => data <= "000000";
				when "001101110010011111" => data <= "000000";
				when "001101111000000000" => data <= "000000";
				when "001101111000000001" => data <= "000000";
				when "001101111000000010" => data <= "000000";
				when "001101111000000011" => data <= "000000";
				when "001101111000000100" => data <= "000000";
				when "001101111000000101" => data <= "000000";
				when "001101111000000110" => data <= "000000";
				when "001101111000000111" => data <= "000000";
				when "001101111000001000" => data <= "000000";
				when "001101111000001001" => data <= "000000";
				when "001101111000001010" => data <= "000000";
				when "001101111000001011" => data <= "000000";
				when "001101111000001100" => data <= "000000";
				when "001101111000001101" => data <= "000000";
				when "001101111000001110" => data <= "000000";
				when "001101111000001111" => data <= "000000";
				when "001101111000010000" => data <= "000000";
				when "001101111000010001" => data <= "000000";
				when "001101111000010010" => data <= "000000";
				when "001101111000010011" => data <= "000000";
				when "001101111000010100" => data <= "000000";
				when "001101111000010101" => data <= "000000";
				when "001101111000010110" => data <= "000000";
				when "001101111000010111" => data <= "000000";
				when "001101111000011000" => data <= "000000";
				when "001101111000011001" => data <= "000000";
				when "001101111000011010" => data <= "000000";
				when "001101111000011011" => data <= "000000";
				when "001101111000011100" => data <= "000000";
				when "001101111000011101" => data <= "000000";
				when "001101111000011110" => data <= "000000";
				when "001101111000011111" => data <= "000000";
				when "001101111000100000" => data <= "000000";
				when "001101111000100001" => data <= "000000";
				when "001101111000100010" => data <= "000000";
				when "001101111000100011" => data <= "000000";
				when "001101111000100100" => data <= "000000";
				when "001101111000100101" => data <= "000000";
				when "001101111000100110" => data <= "000000";
				when "001101111000100111" => data <= "000000";
				when "001101111000101000" => data <= "000000";
				when "001101111000101001" => data <= "000000";
				when "001101111000101010" => data <= "000000";
				when "001101111000101011" => data <= "000000";
				when "001101111000101100" => data <= "000000";
				when "001101111000101101" => data <= "000000";
				when "001101111000101110" => data <= "000000";
				when "001101111000101111" => data <= "000000";
				when "001101111000110000" => data <= "000000";
				when "001101111000110001" => data <= "000000";
				when "001101111000110010" => data <= "000000";
				when "001101111000110011" => data <= "000000";
				when "001101111000110100" => data <= "000000";
				when "001101111000110101" => data <= "000000";
				when "001101111000110110" => data <= "000000";
				when "001101111000110111" => data <= "000000";
				when "001101111000111000" => data <= "000000";
				when "001101111000111001" => data <= "000000";
				when "001101111000111010" => data <= "000000";
				when "001101111000111011" => data <= "000000";
				when "001101111000111100" => data <= "000000";
				when "001101111000111101" => data <= "000000";
				when "001101111000111110" => data <= "000000";
				when "001101111000111111" => data <= "000000";
				when "001101111001000000" => data <= "000000";
				when "001101111001000001" => data <= "000000";
				when "001101111001000010" => data <= "000000";
				when "001101111001000011" => data <= "000000";
				when "001101111001000100" => data <= "000000";
				when "001101111001000101" => data <= "000000";
				when "001101111001000110" => data <= "000000";
				when "001101111001000111" => data <= "000000";
				when "001101111001001000" => data <= "000000";
				when "001101111001001001" => data <= "000000";
				when "001101111001001010" => data <= "000000";
				when "001101111001001011" => data <= "000000";
				when "001101111001001100" => data <= "000000";
				when "001101111001001101" => data <= "000000";
				when "001101111001001110" => data <= "000000";
				when "001101111001001111" => data <= "000000";
				when "001101111001010000" => data <= "000000";
				when "001101111001010001" => data <= "000000";
				when "001101111001010010" => data <= "000000";
				when "001101111001010011" => data <= "000000";
				when "001101111001010100" => data <= "000000";
				when "001101111001010101" => data <= "000000";
				when "001101111001010110" => data <= "000000";
				when "001101111001010111" => data <= "000000";
				when "001101111001011000" => data <= "000000";
				when "001101111001011001" => data <= "000000";
				when "001101111001011010" => data <= "000000";
				when "001101111001011011" => data <= "000000";
				when "001101111001011100" => data <= "000000";
				when "001101111001011101" => data <= "000000";
				when "001101111001011110" => data <= "000000";
				when "001101111001011111" => data <= "000000";
				when "001101111001100000" => data <= "000000";
				when "001101111001100001" => data <= "000000";
				when "001101111001100010" => data <= "000000";
				when "001101111001100011" => data <= "000000";
				when "001101111001100100" => data <= "000000";
				when "001101111001100101" => data <= "000000";
				when "001101111001100110" => data <= "000000";
				when "001101111001100111" => data <= "000000";
				when "001101111001101000" => data <= "000000";
				when "001101111001101001" => data <= "000000";
				when "001101111001101010" => data <= "000000";
				when "001101111001101011" => data <= "000000";
				when "001101111001101100" => data <= "000000";
				when "001101111001101101" => data <= "000000";
				when "001101111001101110" => data <= "000000";
				when "001101111001101111" => data <= "000000";
				when "001101111001110000" => data <= "000000";
				when "001101111001110001" => data <= "000000";
				when "001101111001110010" => data <= "000000";
				when "001101111001110011" => data <= "000000";
				when "001101111001110100" => data <= "000000";
				when "001101111001110101" => data <= "000000";
				when "001101111001110110" => data <= "000000";
				when "001101111001110111" => data <= "000000";
				when "001101111001111000" => data <= "000000";
				when "001101111001111001" => data <= "000000";
				when "001101111001111010" => data <= "000000";
				when "001101111001111011" => data <= "000000";
				when "001101111001111100" => data <= "000000";
				when "001101111001111101" => data <= "000000";
				when "001101111001111110" => data <= "000000";
				when "001101111001111111" => data <= "000000";
				when "001101111010000000" => data <= "000000";
				when "001101111010000001" => data <= "000000";
				when "001101111010000010" => data <= "000000";
				when "001101111010000011" => data <= "000000";
				when "001101111010000100" => data <= "000000";
				when "001101111010000101" => data <= "000000";
				when "001101111010000110" => data <= "000000";
				when "001101111010000111" => data <= "000000";
				when "001101111010001000" => data <= "000000";
				when "001101111010001001" => data <= "000000";
				when "001101111010001010" => data <= "000000";
				when "001101111010001011" => data <= "000000";
				when "001101111010001100" => data <= "000000";
				when "001101111010001101" => data <= "000000";
				when "001101111010001110" => data <= "000000";
				when "001101111010001111" => data <= "000000";
				when "001101111010010000" => data <= "000000";
				when "001101111010010001" => data <= "000000";
				when "001101111010010010" => data <= "000000";
				when "001101111010010011" => data <= "000000";
				when "001101111010010100" => data <= "000000";
				when "001101111010010101" => data <= "000000";
				when "001101111010010110" => data <= "000000";
				when "001101111010010111" => data <= "000000";
				when "001101111010011000" => data <= "000000";
				when "001101111010011001" => data <= "000000";
				when "001101111010011010" => data <= "000000";
				when "001101111010011011" => data <= "000000";
				when "001101111010011100" => data <= "000000";
				when "001101111010011101" => data <= "000000";
				when "001101111010011110" => data <= "000000";
				when "001101111010011111" => data <= "000000";
				when "001110000000000000" => data <= "000000";
				when "001110000000000001" => data <= "000000";
				when "001110000000000010" => data <= "000000";
				when "001110000000000011" => data <= "000000";
				when "001110000000000100" => data <= "000000";
				when "001110000000000101" => data <= "000000";
				when "001110000000000110" => data <= "000000";
				when "001110000000000111" => data <= "000000";
				when "001110000000001000" => data <= "000000";
				when "001110000000001001" => data <= "000000";
				when "001110000000001010" => data <= "000000";
				when "001110000000001011" => data <= "000000";
				when "001110000000001100" => data <= "000000";
				when "001110000000001101" => data <= "000000";
				when "001110000000001110" => data <= "000000";
				when "001110000000001111" => data <= "000000";
				when "001110000000010000" => data <= "000000";
				when "001110000000010001" => data <= "000000";
				when "001110000000010010" => data <= "000000";
				when "001110000000010011" => data <= "000000";
				when "001110000000010100" => data <= "000000";
				when "001110000000010101" => data <= "000000";
				when "001110000000010110" => data <= "000000";
				when "001110000000010111" => data <= "000000";
				when "001110000000011000" => data <= "000000";
				when "001110000000011001" => data <= "000000";
				when "001110000000011010" => data <= "000000";
				when "001110000000011011" => data <= "000000";
				when "001110000000011100" => data <= "000000";
				when "001110000000011101" => data <= "000000";
				when "001110000000011110" => data <= "000000";
				when "001110000000011111" => data <= "000000";
				when "001110000000100000" => data <= "000000";
				when "001110000000100001" => data <= "000000";
				when "001110000000100010" => data <= "000000";
				when "001110000000100011" => data <= "000000";
				when "001110000000100100" => data <= "000000";
				when "001110000000100101" => data <= "000000";
				when "001110000000100110" => data <= "000000";
				when "001110000000100111" => data <= "000000";
				when "001110000000101000" => data <= "000000";
				when "001110000000101001" => data <= "000000";
				when "001110000000101010" => data <= "000000";
				when "001110000000101011" => data <= "000000";
				when "001110000000101100" => data <= "000000";
				when "001110000000101101" => data <= "000000";
				when "001110000000101110" => data <= "000000";
				when "001110000000101111" => data <= "000000";
				when "001110000000110000" => data <= "000000";
				when "001110000000110001" => data <= "000000";
				when "001110000000110010" => data <= "000000";
				when "001110000000110011" => data <= "000000";
				when "001110000000110100" => data <= "000000";
				when "001110000000110101" => data <= "000000";
				when "001110000000110110" => data <= "000000";
				when "001110000000110111" => data <= "000000";
				when "001110000000111000" => data <= "000000";
				when "001110000000111001" => data <= "000000";
				when "001110000000111010" => data <= "000000";
				when "001110000000111011" => data <= "000000";
				when "001110000000111100" => data <= "000000";
				when "001110000000111101" => data <= "000000";
				when "001110000000111110" => data <= "000000";
				when "001110000000111111" => data <= "000000";
				when "001110000001000000" => data <= "000000";
				when "001110000001000001" => data <= "000000";
				when "001110000001000010" => data <= "000000";
				when "001110000001000011" => data <= "000000";
				when "001110000001000100" => data <= "000000";
				when "001110000001000101" => data <= "000000";
				when "001110000001000110" => data <= "000000";
				when "001110000001000111" => data <= "000000";
				when "001110000001001000" => data <= "000000";
				when "001110000001001001" => data <= "000000";
				when "001110000001001010" => data <= "000000";
				when "001110000001001011" => data <= "000000";
				when "001110000001001100" => data <= "000000";
				when "001110000001001101" => data <= "000000";
				when "001110000001001110" => data <= "000000";
				when "001110000001001111" => data <= "000000";
				when "001110000001010000" => data <= "000000";
				when "001110000001010001" => data <= "000000";
				when "001110000001010010" => data <= "000000";
				when "001110000001010011" => data <= "000000";
				when "001110000001010100" => data <= "000000";
				when "001110000001010101" => data <= "000000";
				when "001110000001010110" => data <= "000000";
				when "001110000001010111" => data <= "000000";
				when "001110000001011000" => data <= "000000";
				when "001110000001011001" => data <= "000000";
				when "001110000001011010" => data <= "000000";
				when "001110000001011011" => data <= "000000";
				when "001110000001011100" => data <= "000000";
				when "001110000001011101" => data <= "000000";
				when "001110000001011110" => data <= "000000";
				when "001110000001011111" => data <= "000000";
				when "001110000001100000" => data <= "000000";
				when "001110000001100001" => data <= "000000";
				when "001110000001100010" => data <= "000000";
				when "001110000001100011" => data <= "000000";
				when "001110000001100100" => data <= "000000";
				when "001110000001100101" => data <= "000000";
				when "001110000001100110" => data <= "000000";
				when "001110000001100111" => data <= "000000";
				when "001110000001101000" => data <= "000000";
				when "001110000001101001" => data <= "000000";
				when "001110000001101010" => data <= "000000";
				when "001110000001101011" => data <= "000000";
				when "001110000001101100" => data <= "000000";
				when "001110000001101101" => data <= "000000";
				when "001110000001101110" => data <= "000000";
				when "001110000001101111" => data <= "000000";
				when "001110000001110000" => data <= "000000";
				when "001110000001110001" => data <= "000000";
				when "001110000001110010" => data <= "000000";
				when "001110000001110011" => data <= "000000";
				when "001110000001110100" => data <= "000000";
				when "001110000001110101" => data <= "000000";
				when "001110000001110110" => data <= "000000";
				when "001110000001110111" => data <= "000000";
				when "001110000001111000" => data <= "000000";
				when "001110000001111001" => data <= "000000";
				when "001110000001111010" => data <= "000000";
				when "001110000001111011" => data <= "000000";
				when "001110000001111100" => data <= "000000";
				when "001110000001111101" => data <= "000000";
				when "001110000001111110" => data <= "000000";
				when "001110000001111111" => data <= "000000";
				when "001110000010000000" => data <= "000000";
				when "001110000010000001" => data <= "000000";
				when "001110000010000010" => data <= "000000";
				when "001110000010000011" => data <= "000000";
				when "001110000010000100" => data <= "000000";
				when "001110000010000101" => data <= "000000";
				when "001110000010000110" => data <= "000000";
				when "001110000010000111" => data <= "000000";
				when "001110000010001000" => data <= "000000";
				when "001110000010001001" => data <= "000000";
				when "001110000010001010" => data <= "000000";
				when "001110000010001011" => data <= "000000";
				when "001110000010001100" => data <= "000000";
				when "001110000010001101" => data <= "000000";
				when "001110000010001110" => data <= "000000";
				when "001110000010001111" => data <= "000000";
				when "001110000010010000" => data <= "000000";
				when "001110000010010001" => data <= "000000";
				when "001110000010010010" => data <= "000000";
				when "001110000010010011" => data <= "000000";
				when "001110000010010100" => data <= "000000";
				when "001110000010010101" => data <= "000000";
				when "001110000010010110" => data <= "000000";
				when "001110000010010111" => data <= "000000";
				when "001110000010011000" => data <= "000000";
				when "001110000010011001" => data <= "000000";
				when "001110000010011010" => data <= "000000";
				when "001110000010011011" => data <= "000000";
				when "001110000010011100" => data <= "000000";
				when "001110000010011101" => data <= "000000";
				when "001110000010011110" => data <= "000000";
				when "001110000010011111" => data <= "000000";
				when "001110001000000000" => data <= "000000";
				when "001110001000000001" => data <= "000000";
				when "001110001000000010" => data <= "000000";
				when "001110001000000011" => data <= "000000";
				when "001110001000000100" => data <= "000000";
				when "001110001000000101" => data <= "000000";
				when "001110001000000110" => data <= "000000";
				when "001110001000000111" => data <= "000000";
				when "001110001000001000" => data <= "000000";
				when "001110001000001001" => data <= "000000";
				when "001110001000001010" => data <= "000000";
				when "001110001000001011" => data <= "000000";
				when "001110001000001100" => data <= "000000";
				when "001110001000001101" => data <= "000000";
				when "001110001000001110" => data <= "000000";
				when "001110001000001111" => data <= "000000";
				when "001110001000010000" => data <= "000000";
				when "001110001000010001" => data <= "000000";
				when "001110001000010010" => data <= "000000";
				when "001110001000010011" => data <= "000000";
				when "001110001000010100" => data <= "000000";
				when "001110001000010101" => data <= "000000";
				when "001110001000010110" => data <= "000000";
				when "001110001000010111" => data <= "000000";
				when "001110001000011000" => data <= "000000";
				when "001110001000011001" => data <= "000000";
				when "001110001000011010" => data <= "000000";
				when "001110001000011011" => data <= "000000";
				when "001110001000011100" => data <= "000000";
				when "001110001000011101" => data <= "000000";
				when "001110001000011110" => data <= "000000";
				when "001110001000011111" => data <= "000000";
				when "001110001000100000" => data <= "000000";
				when "001110001000100001" => data <= "000000";
				when "001110001000100010" => data <= "000000";
				when "001110001000100011" => data <= "000000";
				when "001110001000100100" => data <= "000000";
				when "001110001000100101" => data <= "000000";
				when "001110001000100110" => data <= "000000";
				when "001110001000100111" => data <= "000000";
				when "001110001000101000" => data <= "000000";
				when "001110001000101001" => data <= "000000";
				when "001110001000101010" => data <= "000000";
				when "001110001000101011" => data <= "000000";
				when "001110001000101100" => data <= "000000";
				when "001110001000101101" => data <= "000000";
				when "001110001000101110" => data <= "000000";
				when "001110001000101111" => data <= "000000";
				when "001110001000110000" => data <= "000000";
				when "001110001000110001" => data <= "000000";
				when "001110001000110010" => data <= "000000";
				when "001110001000110011" => data <= "000000";
				when "001110001000110100" => data <= "000000";
				when "001110001000110101" => data <= "000000";
				when "001110001000110110" => data <= "000000";
				when "001110001000110111" => data <= "000000";
				when "001110001000111000" => data <= "000000";
				when "001110001000111001" => data <= "000000";
				when "001110001000111010" => data <= "000000";
				when "001110001000111011" => data <= "000000";
				when "001110001000111100" => data <= "000000";
				when "001110001000111101" => data <= "000000";
				when "001110001000111110" => data <= "000000";
				when "001110001000111111" => data <= "000000";
				when "001110001001000000" => data <= "000000";
				when "001110001001000001" => data <= "000000";
				when "001110001001000010" => data <= "000000";
				when "001110001001000011" => data <= "000000";
				when "001110001001000100" => data <= "000000";
				when "001110001001000101" => data <= "000000";
				when "001110001001000110" => data <= "000000";
				when "001110001001000111" => data <= "000000";
				when "001110001001001000" => data <= "000000";
				when "001110001001001001" => data <= "000000";
				when "001110001001001010" => data <= "000000";
				when "001110001001001011" => data <= "000000";
				when "001110001001001100" => data <= "000000";
				when "001110001001001101" => data <= "000000";
				when "001110001001001110" => data <= "000000";
				when "001110001001001111" => data <= "000000";
				when "001110001001010000" => data <= "000000";
				when "001110001001010001" => data <= "000000";
				when "001110001001010010" => data <= "000000";
				when "001110001001010011" => data <= "000000";
				when "001110001001010100" => data <= "000000";
				when "001110001001010101" => data <= "000000";
				when "001110001001010110" => data <= "000000";
				when "001110001001010111" => data <= "000000";
				when "001110001001011000" => data <= "000000";
				when "001110001001011001" => data <= "000000";
				when "001110001001011010" => data <= "000000";
				when "001110001001011011" => data <= "000000";
				when "001110001001011100" => data <= "000000";
				when "001110001001011101" => data <= "000000";
				when "001110001001011110" => data <= "000000";
				when "001110001001011111" => data <= "000000";
				when "001110001001100000" => data <= "000000";
				when "001110001001100001" => data <= "000000";
				when "001110001001100010" => data <= "000000";
				when "001110001001100011" => data <= "000000";
				when "001110001001100100" => data <= "000000";
				when "001110001001100101" => data <= "000000";
				when "001110001001100110" => data <= "000000";
				when "001110001001100111" => data <= "000000";
				when "001110001001101000" => data <= "000000";
				when "001110001001101001" => data <= "000000";
				when "001110001001101010" => data <= "000000";
				when "001110001001101011" => data <= "000000";
				when "001110001001101100" => data <= "000000";
				when "001110001001101101" => data <= "000000";
				when "001110001001101110" => data <= "000000";
				when "001110001001101111" => data <= "000000";
				when "001110001001110000" => data <= "000000";
				when "001110001001110001" => data <= "000000";
				when "001110001001110010" => data <= "000000";
				when "001110001001110011" => data <= "000000";
				when "001110001001110100" => data <= "000000";
				when "001110001001110101" => data <= "000000";
				when "001110001001110110" => data <= "000000";
				when "001110001001110111" => data <= "000000";
				when "001110001001111000" => data <= "000000";
				when "001110001001111001" => data <= "000000";
				when "001110001001111010" => data <= "000000";
				when "001110001001111011" => data <= "000000";
				when "001110001001111100" => data <= "000000";
				when "001110001001111101" => data <= "000000";
				when "001110001001111110" => data <= "000000";
				when "001110001001111111" => data <= "000000";
				when "001110001010000000" => data <= "000000";
				when "001110001010000001" => data <= "000000";
				when "001110001010000010" => data <= "000000";
				when "001110001010000011" => data <= "000000";
				when "001110001010000100" => data <= "000000";
				when "001110001010000101" => data <= "000000";
				when "001110001010000110" => data <= "000000";
				when "001110001010000111" => data <= "000000";
				when "001110001010001000" => data <= "000000";
				when "001110001010001001" => data <= "000000";
				when "001110001010001010" => data <= "000000";
				when "001110001010001011" => data <= "000000";
				when "001110001010001100" => data <= "000000";
				when "001110001010001101" => data <= "000000";
				when "001110001010001110" => data <= "000000";
				when "001110001010001111" => data <= "000000";
				when "001110001010010000" => data <= "000000";
				when "001110001010010001" => data <= "000000";
				when "001110001010010010" => data <= "000000";
				when "001110001010010011" => data <= "000000";
				when "001110001010010100" => data <= "000000";
				when "001110001010010101" => data <= "000000";
				when "001110001010010110" => data <= "000000";
				when "001110001010010111" => data <= "000000";
				when "001110001010011000" => data <= "000000";
				when "001110001010011001" => data <= "000000";
				when "001110001010011010" => data <= "000000";
				when "001110001010011011" => data <= "000000";
				when "001110001010011100" => data <= "000000";
				when "001110001010011101" => data <= "000000";
				when "001110001010011110" => data <= "000000";
				when "001110001010011111" => data <= "000000";
				when "001110010000000000" => data <= "000000";
				when "001110010000000001" => data <= "000000";
				when "001110010000000010" => data <= "000000";
				when "001110010000000011" => data <= "000000";
				when "001110010000000100" => data <= "000000";
				when "001110010000000101" => data <= "000000";
				when "001110010000000110" => data <= "000000";
				when "001110010000000111" => data <= "000000";
				when "001110010000001000" => data <= "000000";
				when "001110010000001001" => data <= "000000";
				when "001110010000001010" => data <= "000000";
				when "001110010000001011" => data <= "000000";
				when "001110010000001100" => data <= "000000";
				when "001110010000001101" => data <= "000000";
				when "001110010000001110" => data <= "000000";
				when "001110010000001111" => data <= "000000";
				when "001110010000010000" => data <= "000000";
				when "001110010000010001" => data <= "000000";
				when "001110010000010010" => data <= "000000";
				when "001110010000010011" => data <= "000000";
				when "001110010000010100" => data <= "000000";
				when "001110010000010101" => data <= "000000";
				when "001110010000010110" => data <= "000000";
				when "001110010000010111" => data <= "000000";
				when "001110010000011000" => data <= "000000";
				when "001110010000011001" => data <= "000000";
				when "001110010000011010" => data <= "000000";
				when "001110010000011011" => data <= "000000";
				when "001110010000011100" => data <= "000000";
				when "001110010000011101" => data <= "000000";
				when "001110010000011110" => data <= "000000";
				when "001110010000011111" => data <= "000000";
				when "001110010000100000" => data <= "000000";
				when "001110010000100001" => data <= "000000";
				when "001110010000100010" => data <= "000000";
				when "001110010000100011" => data <= "000000";
				when "001110010000100100" => data <= "000000";
				when "001110010000100101" => data <= "000000";
				when "001110010000100110" => data <= "000000";
				when "001110010000100111" => data <= "000000";
				when "001110010000101000" => data <= "000000";
				when "001110010000101001" => data <= "000000";
				when "001110010000101010" => data <= "000000";
				when "001110010000101011" => data <= "000000";
				when "001110010000101100" => data <= "000000";
				when "001110010000101101" => data <= "000000";
				when "001110010000101110" => data <= "000000";
				when "001110010000101111" => data <= "000000";
				when "001110010000110000" => data <= "000000";
				when "001110010000110001" => data <= "000000";
				when "001110010000110010" => data <= "000000";
				when "001110010000110011" => data <= "000000";
				when "001110010000110100" => data <= "000000";
				when "001110010000110101" => data <= "000000";
				when "001110010000110110" => data <= "000000";
				when "001110010000110111" => data <= "000000";
				when "001110010000111000" => data <= "000000";
				when "001110010000111001" => data <= "000000";
				when "001110010000111010" => data <= "000000";
				when "001110010000111011" => data <= "000000";
				when "001110010000111100" => data <= "000000";
				when "001110010000111101" => data <= "000000";
				when "001110010000111110" => data <= "000000";
				when "001110010000111111" => data <= "000000";
				when "001110010001000000" => data <= "000000";
				when "001110010001000001" => data <= "000000";
				when "001110010001000010" => data <= "000000";
				when "001110010001000011" => data <= "000000";
				when "001110010001000100" => data <= "000000";
				when "001110010001000101" => data <= "000000";
				when "001110010001000110" => data <= "000000";
				when "001110010001000111" => data <= "000000";
				when "001110010001001000" => data <= "000000";
				when "001110010001001001" => data <= "000000";
				when "001110010001001010" => data <= "000000";
				when "001110010001001011" => data <= "000000";
				when "001110010001001100" => data <= "000000";
				when "001110010001001101" => data <= "000000";
				when "001110010001001110" => data <= "000000";
				when "001110010001001111" => data <= "000000";
				when "001110010001010000" => data <= "000000";
				when "001110010001010001" => data <= "000000";
				when "001110010001010010" => data <= "000000";
				when "001110010001010011" => data <= "000000";
				when "001110010001010100" => data <= "000000";
				when "001110010001010101" => data <= "000000";
				when "001110010001010110" => data <= "000000";
				when "001110010001010111" => data <= "000000";
				when "001110010001011000" => data <= "000000";
				when "001110010001011001" => data <= "000000";
				when "001110010001011010" => data <= "000000";
				when "001110010001011011" => data <= "000000";
				when "001110010001011100" => data <= "000000";
				when "001110010001011101" => data <= "000000";
				when "001110010001011110" => data <= "000000";
				when "001110010001011111" => data <= "000000";
				when "001110010001100000" => data <= "000000";
				when "001110010001100001" => data <= "000000";
				when "001110010001100010" => data <= "000000";
				when "001110010001100011" => data <= "000000";
				when "001110010001100100" => data <= "000000";
				when "001110010001100101" => data <= "000000";
				when "001110010001100110" => data <= "000000";
				when "001110010001100111" => data <= "000000";
				when "001110010001101000" => data <= "000000";
				when "001110010001101001" => data <= "000000";
				when "001110010001101010" => data <= "000000";
				when "001110010001101011" => data <= "000000";
				when "001110010001101100" => data <= "000000";
				when "001110010001101101" => data <= "000000";
				when "001110010001101110" => data <= "000000";
				when "001110010001101111" => data <= "000000";
				when "001110010001110000" => data <= "000000";
				when "001110010001110001" => data <= "000000";
				when "001110010001110010" => data <= "000000";
				when "001110010001110011" => data <= "000000";
				when "001110010001110100" => data <= "000000";
				when "001110010001110101" => data <= "000000";
				when "001110010001110110" => data <= "000000";
				when "001110010001110111" => data <= "000000";
				when "001110010001111000" => data <= "000000";
				when "001110010001111001" => data <= "000000";
				when "001110010001111010" => data <= "000000";
				when "001110010001111011" => data <= "000000";
				when "001110010001111100" => data <= "000000";
				when "001110010001111101" => data <= "000000";
				when "001110010001111110" => data <= "000000";
				when "001110010001111111" => data <= "000000";
				when "001110010010000000" => data <= "000000";
				when "001110010010000001" => data <= "000000";
				when "001110010010000010" => data <= "000000";
				when "001110010010000011" => data <= "000000";
				when "001110010010000100" => data <= "000000";
				when "001110010010000101" => data <= "000000";
				when "001110010010000110" => data <= "000000";
				when "001110010010000111" => data <= "000000";
				when "001110010010001000" => data <= "000000";
				when "001110010010001001" => data <= "000000";
				when "001110010010001010" => data <= "000000";
				when "001110010010001011" => data <= "000000";
				when "001110010010001100" => data <= "000000";
				when "001110010010001101" => data <= "000000";
				when "001110010010001110" => data <= "000000";
				when "001110010010001111" => data <= "000000";
				when "001110010010010000" => data <= "000000";
				when "001110010010010001" => data <= "000000";
				when "001110010010010010" => data <= "000000";
				when "001110010010010011" => data <= "000000";
				when "001110010010010100" => data <= "000000";
				when "001110010010010101" => data <= "000000";
				when "001110010010010110" => data <= "000000";
				when "001110010010010111" => data <= "000000";
				when "001110010010011000" => data <= "000000";
				when "001110010010011001" => data <= "000000";
				when "001110010010011010" => data <= "000000";
				when "001110010010011011" => data <= "000000";
				when "001110010010011100" => data <= "000000";
				when "001110010010011101" => data <= "000000";
				when "001110010010011110" => data <= "000000";
				when "001110010010011111" => data <= "000000";
				when "001110011000000000" => data <= "000000";
				when "001110011000000001" => data <= "000000";
				when "001110011000000010" => data <= "000000";
				when "001110011000000011" => data <= "000000";
				when "001110011000000100" => data <= "000000";
				when "001110011000000101" => data <= "000000";
				when "001110011000000110" => data <= "000000";
				when "001110011000000111" => data <= "000000";
				when "001110011000001000" => data <= "000000";
				when "001110011000001001" => data <= "000000";
				when "001110011000001010" => data <= "000000";
				when "001110011000001011" => data <= "000000";
				when "001110011000001100" => data <= "000000";
				when "001110011000001101" => data <= "000000";
				when "001110011000001110" => data <= "000000";
				when "001110011000001111" => data <= "000000";
				when "001110011000010000" => data <= "000000";
				when "001110011000010001" => data <= "000000";
				when "001110011000010010" => data <= "000000";
				when "001110011000010011" => data <= "000000";
				when "001110011000010100" => data <= "000000";
				when "001110011000010101" => data <= "000000";
				when "001110011000010110" => data <= "000000";
				when "001110011000010111" => data <= "000000";
				when "001110011000011000" => data <= "000000";
				when "001110011000011001" => data <= "000000";
				when "001110011000011010" => data <= "000000";
				when "001110011000011011" => data <= "000000";
				when "001110011000011100" => data <= "000000";
				when "001110011000011101" => data <= "000000";
				when "001110011000011110" => data <= "000000";
				when "001110011000011111" => data <= "000000";
				when "001110011000100000" => data <= "000000";
				when "001110011000100001" => data <= "000000";
				when "001110011000100010" => data <= "000000";
				when "001110011000100011" => data <= "000000";
				when "001110011000100100" => data <= "000000";
				when "001110011000100101" => data <= "000000";
				when "001110011000100110" => data <= "000000";
				when "001110011000100111" => data <= "000000";
				when "001110011000101000" => data <= "000000";
				when "001110011000101001" => data <= "000000";
				when "001110011000101010" => data <= "000000";
				when "001110011000101011" => data <= "000000";
				when "001110011000101100" => data <= "000000";
				when "001110011000101101" => data <= "000000";
				when "001110011000101110" => data <= "000000";
				when "001110011000101111" => data <= "000000";
				when "001110011000110000" => data <= "000000";
				when "001110011000110001" => data <= "000000";
				when "001110011000110010" => data <= "000000";
				when "001110011000110011" => data <= "000000";
				when "001110011000110100" => data <= "000000";
				when "001110011000110101" => data <= "000000";
				when "001110011000110110" => data <= "000000";
				when "001110011000110111" => data <= "000000";
				when "001110011000111000" => data <= "000000";
				when "001110011000111001" => data <= "000000";
				when "001110011000111010" => data <= "000000";
				when "001110011000111011" => data <= "000000";
				when "001110011000111100" => data <= "000000";
				when "001110011000111101" => data <= "000000";
				when "001110011000111110" => data <= "000000";
				when "001110011000111111" => data <= "000000";
				when "001110011001000000" => data <= "000000";
				when "001110011001000001" => data <= "000000";
				when "001110011001000010" => data <= "000000";
				when "001110011001000011" => data <= "000000";
				when "001110011001000100" => data <= "000000";
				when "001110011001000101" => data <= "000000";
				when "001110011001000110" => data <= "000000";
				when "001110011001000111" => data <= "000000";
				when "001110011001001000" => data <= "000000";
				when "001110011001001001" => data <= "000000";
				when "001110011001001010" => data <= "000000";
				when "001110011001001011" => data <= "000000";
				when "001110011001001100" => data <= "000000";
				when "001110011001001101" => data <= "000000";
				when "001110011001001110" => data <= "000000";
				when "001110011001001111" => data <= "000000";
				when "001110011001010000" => data <= "000000";
				when "001110011001010001" => data <= "000000";
				when "001110011001010010" => data <= "000000";
				when "001110011001010011" => data <= "000000";
				when "001110011001010100" => data <= "000000";
				when "001110011001010101" => data <= "000000";
				when "001110011001010110" => data <= "000000";
				when "001110011001010111" => data <= "000000";
				when "001110011001011000" => data <= "000000";
				when "001110011001011001" => data <= "000000";
				when "001110011001011010" => data <= "000000";
				when "001110011001011011" => data <= "000000";
				when "001110011001011100" => data <= "000000";
				when "001110011001011101" => data <= "000000";
				when "001110011001011110" => data <= "000000";
				when "001110011001011111" => data <= "000000";
				when "001110011001100000" => data <= "000000";
				when "001110011001100001" => data <= "000000";
				when "001110011001100010" => data <= "000000";
				when "001110011001100011" => data <= "000000";
				when "001110011001100100" => data <= "000000";
				when "001110011001100101" => data <= "000000";
				when "001110011001100110" => data <= "000000";
				when "001110011001100111" => data <= "000000";
				when "001110011001101000" => data <= "000000";
				when "001110011001101001" => data <= "000000";
				when "001110011001101010" => data <= "000000";
				when "001110011001101011" => data <= "000000";
				when "001110011001101100" => data <= "000000";
				when "001110011001101101" => data <= "000000";
				when "001110011001101110" => data <= "000000";
				when "001110011001101111" => data <= "000000";
				when "001110011001110000" => data <= "000000";
				when "001110011001110001" => data <= "000000";
				when "001110011001110010" => data <= "000000";
				when "001110011001110011" => data <= "000000";
				when "001110011001110100" => data <= "000000";
				when "001110011001110101" => data <= "000000";
				when "001110011001110110" => data <= "000000";
				when "001110011001110111" => data <= "000000";
				when "001110011001111000" => data <= "000000";
				when "001110011001111001" => data <= "000000";
				when "001110011001111010" => data <= "000000";
				when "001110011001111011" => data <= "000000";
				when "001110011001111100" => data <= "000000";
				when "001110011001111101" => data <= "000000";
				when "001110011001111110" => data <= "000000";
				when "001110011001111111" => data <= "000000";
				when "001110011010000000" => data <= "000000";
				when "001110011010000001" => data <= "000000";
				when "001110011010000010" => data <= "000000";
				when "001110011010000011" => data <= "000000";
				when "001110011010000100" => data <= "000000";
				when "001110011010000101" => data <= "000000";
				when "001110011010000110" => data <= "000000";
				when "001110011010000111" => data <= "000000";
				when "001110011010001000" => data <= "000000";
				when "001110011010001001" => data <= "000000";
				when "001110011010001010" => data <= "000000";
				when "001110011010001011" => data <= "000000";
				when "001110011010001100" => data <= "000000";
				when "001110011010001101" => data <= "000000";
				when "001110011010001110" => data <= "000000";
				when "001110011010001111" => data <= "000000";
				when "001110011010010000" => data <= "000000";
				when "001110011010010001" => data <= "000000";
				when "001110011010010010" => data <= "000000";
				when "001110011010010011" => data <= "000000";
				when "001110011010010100" => data <= "000000";
				when "001110011010010101" => data <= "000000";
				when "001110011010010110" => data <= "000000";
				when "001110011010010111" => data <= "000000";
				when "001110011010011000" => data <= "000000";
				when "001110011010011001" => data <= "000000";
				when "001110011010011010" => data <= "000000";
				when "001110011010011011" => data <= "000000";
				when "001110011010011100" => data <= "000000";
				when "001110011010011101" => data <= "000000";
				when "001110011010011110" => data <= "000000";
				when "001110011010011111" => data <= "000000";
				when "001110100000000000" => data <= "000000";
				when "001110100000000001" => data <= "000000";
				when "001110100000000010" => data <= "000000";
				when "001110100000000011" => data <= "000000";
				when "001110100000000100" => data <= "000000";
				when "001110100000000101" => data <= "000000";
				when "001110100000000110" => data <= "000000";
				when "001110100000000111" => data <= "000000";
				when "001110100000001000" => data <= "000000";
				when "001110100000001001" => data <= "000000";
				when "001110100000001010" => data <= "000000";
				when "001110100000001011" => data <= "000000";
				when "001110100000001100" => data <= "000000";
				when "001110100000001101" => data <= "000000";
				when "001110100000001110" => data <= "000000";
				when "001110100000001111" => data <= "000000";
				when "001110100000010000" => data <= "000000";
				when "001110100000010001" => data <= "000000";
				when "001110100000010010" => data <= "000000";
				when "001110100000010011" => data <= "000000";
				when "001110100000010100" => data <= "000000";
				when "001110100000010101" => data <= "000000";
				when "001110100000010110" => data <= "000000";
				when "001110100000010111" => data <= "000000";
				when "001110100000011000" => data <= "000000";
				when "001110100000011001" => data <= "000000";
				when "001110100000011010" => data <= "000000";
				when "001110100000011011" => data <= "000000";
				when "001110100000011100" => data <= "000000";
				when "001110100000011101" => data <= "000000";
				when "001110100000011110" => data <= "000000";
				when "001110100000011111" => data <= "000000";
				when "001110100000100000" => data <= "000000";
				when "001110100000100001" => data <= "000000";
				when "001110100000100010" => data <= "000000";
				when "001110100000100011" => data <= "000000";
				when "001110100000100100" => data <= "000000";
				when "001110100000100101" => data <= "000000";
				when "001110100000100110" => data <= "000000";
				when "001110100000100111" => data <= "000000";
				when "001110100000101000" => data <= "000000";
				when "001110100000101001" => data <= "000000";
				when "001110100000101010" => data <= "000000";
				when "001110100000101011" => data <= "000000";
				when "001110100000101100" => data <= "000000";
				when "001110100000101101" => data <= "000000";
				when "001110100000101110" => data <= "000000";
				when "001110100000101111" => data <= "000000";
				when "001110100000110000" => data <= "000000";
				when "001110100000110001" => data <= "000000";
				when "001110100000110010" => data <= "000000";
				when "001110100000110011" => data <= "000000";
				when "001110100000110100" => data <= "000000";
				when "001110100000110101" => data <= "000000";
				when "001110100000110110" => data <= "000000";
				when "001110100000110111" => data <= "000000";
				when "001110100000111000" => data <= "000000";
				when "001110100000111001" => data <= "000000";
				when "001110100000111010" => data <= "000000";
				when "001110100000111011" => data <= "000000";
				when "001110100000111100" => data <= "000000";
				when "001110100000111101" => data <= "000000";
				when "001110100000111110" => data <= "000000";
				when "001110100000111111" => data <= "000000";
				when "001110100001000000" => data <= "000000";
				when "001110100001000001" => data <= "000000";
				when "001110100001000010" => data <= "000000";
				when "001110100001000011" => data <= "000000";
				when "001110100001000100" => data <= "000000";
				when "001110100001000101" => data <= "000000";
				when "001110100001000110" => data <= "000000";
				when "001110100001000111" => data <= "000000";
				when "001110100001001000" => data <= "000000";
				when "001110100001001001" => data <= "000000";
				when "001110100001001010" => data <= "000000";
				when "001110100001001011" => data <= "000000";
				when "001110100001001100" => data <= "000000";
				when "001110100001001101" => data <= "000000";
				when "001110100001001110" => data <= "000000";
				when "001110100001001111" => data <= "000000";
				when "001110100001010000" => data <= "000000";
				when "001110100001010001" => data <= "000000";
				when "001110100001010010" => data <= "000000";
				when "001110100001010011" => data <= "000000";
				when "001110100001010100" => data <= "000000";
				when "001110100001010101" => data <= "000000";
				when "001110100001010110" => data <= "000000";
				when "001110100001010111" => data <= "000000";
				when "001110100001011000" => data <= "000000";
				when "001110100001011001" => data <= "000000";
				when "001110100001011010" => data <= "000000";
				when "001110100001011011" => data <= "000000";
				when "001110100001011100" => data <= "000000";
				when "001110100001011101" => data <= "000000";
				when "001110100001011110" => data <= "000000";
				when "001110100001011111" => data <= "000000";
				when "001110100001100000" => data <= "000000";
				when "001110100001100001" => data <= "000000";
				when "001110100001100010" => data <= "000000";
				when "001110100001100011" => data <= "000000";
				when "001110100001100100" => data <= "000000";
				when "001110100001100101" => data <= "000000";
				when "001110100001100110" => data <= "000000";
				when "001110100001100111" => data <= "000000";
				when "001110100001101000" => data <= "000000";
				when "001110100001101001" => data <= "000000";
				when "001110100001101010" => data <= "000000";
				when "001110100001101011" => data <= "000000";
				when "001110100001101100" => data <= "000000";
				when "001110100001101101" => data <= "000000";
				when "001110100001101110" => data <= "000000";
				when "001110100001101111" => data <= "000000";
				when "001110100001110000" => data <= "000000";
				when "001110100001110001" => data <= "000000";
				when "001110100001110010" => data <= "000000";
				when "001110100001110011" => data <= "000000";
				when "001110100001110100" => data <= "000000";
				when "001110100001110101" => data <= "000000";
				when "001110100001110110" => data <= "000000";
				when "001110100001110111" => data <= "000000";
				when "001110100001111000" => data <= "000000";
				when "001110100001111001" => data <= "000000";
				when "001110100001111010" => data <= "000000";
				when "001110100001111011" => data <= "000000";
				when "001110100001111100" => data <= "000000";
				when "001110100001111101" => data <= "000000";
				when "001110100001111110" => data <= "000000";
				when "001110100001111111" => data <= "000000";
				when "001110100010000000" => data <= "000000";
				when "001110100010000001" => data <= "000000";
				when "001110100010000010" => data <= "000000";
				when "001110100010000011" => data <= "000000";
				when "001110100010000100" => data <= "000000";
				when "001110100010000101" => data <= "000000";
				when "001110100010000110" => data <= "000000";
				when "001110100010000111" => data <= "000000";
				when "001110100010001000" => data <= "000000";
				when "001110100010001001" => data <= "000000";
				when "001110100010001010" => data <= "000000";
				when "001110100010001011" => data <= "000000";
				when "001110100010001100" => data <= "000000";
				when "001110100010001101" => data <= "000000";
				when "001110100010001110" => data <= "000000";
				when "001110100010001111" => data <= "000000";
				when "001110100010010000" => data <= "000000";
				when "001110100010010001" => data <= "000000";
				when "001110100010010010" => data <= "000000";
				when "001110100010010011" => data <= "000000";
				when "001110100010010100" => data <= "000000";
				when "001110100010010101" => data <= "000000";
				when "001110100010010110" => data <= "000000";
				when "001110100010010111" => data <= "000000";
				when "001110100010011000" => data <= "000000";
				when "001110100010011001" => data <= "000000";
				when "001110100010011010" => data <= "000000";
				when "001110100010011011" => data <= "000000";
				when "001110100010011100" => data <= "000000";
				when "001110100010011101" => data <= "000000";
				when "001110100010011110" => data <= "000000";
				when "001110100010011111" => data <= "000000";
				when "001110101000000000" => data <= "000000";
				when "001110101000000001" => data <= "000000";
				when "001110101000000010" => data <= "000000";
				when "001110101000000011" => data <= "000000";
				when "001110101000000100" => data <= "000000";
				when "001110101000000101" => data <= "000000";
				when "001110101000000110" => data <= "000000";
				when "001110101000000111" => data <= "000000";
				when "001110101000001000" => data <= "000000";
				when "001110101000001001" => data <= "000000";
				when "001110101000001010" => data <= "000000";
				when "001110101000001011" => data <= "000000";
				when "001110101000001100" => data <= "000000";
				when "001110101000001101" => data <= "000000";
				when "001110101000001110" => data <= "000000";
				when "001110101000001111" => data <= "000000";
				when "001110101000010000" => data <= "000000";
				when "001110101000010001" => data <= "000000";
				when "001110101000010010" => data <= "000000";
				when "001110101000010011" => data <= "000000";
				when "001110101000010100" => data <= "000000";
				when "001110101000010101" => data <= "000000";
				when "001110101000010110" => data <= "000000";
				when "001110101000010111" => data <= "000000";
				when "001110101000011000" => data <= "000000";
				when "001110101000011001" => data <= "000000";
				when "001110101000011010" => data <= "000000";
				when "001110101000011011" => data <= "000000";
				when "001110101000011100" => data <= "000000";
				when "001110101000011101" => data <= "000000";
				when "001110101000011110" => data <= "000000";
				when "001110101000011111" => data <= "000000";
				when "001110101000100000" => data <= "000000";
				when "001110101000100001" => data <= "000000";
				when "001110101000100010" => data <= "000000";
				when "001110101000100011" => data <= "000000";
				when "001110101000100100" => data <= "000000";
				when "001110101000100101" => data <= "000000";
				when "001110101000100110" => data <= "000000";
				when "001110101000100111" => data <= "000000";
				when "001110101000101000" => data <= "000000";
				when "001110101000101001" => data <= "000000";
				when "001110101000101010" => data <= "000000";
				when "001110101000101011" => data <= "000000";
				when "001110101000101100" => data <= "000000";
				when "001110101000101101" => data <= "000000";
				when "001110101000101110" => data <= "000000";
				when "001110101000101111" => data <= "000000";
				when "001110101000110000" => data <= "000000";
				when "001110101000110001" => data <= "000000";
				when "001110101000110010" => data <= "000000";
				when "001110101000110011" => data <= "000000";
				when "001110101000110100" => data <= "000000";
				when "001110101000110101" => data <= "000000";
				when "001110101000110110" => data <= "000000";
				when "001110101000110111" => data <= "000000";
				when "001110101000111000" => data <= "000000";
				when "001110101000111001" => data <= "000000";
				when "001110101000111010" => data <= "000000";
				when "001110101000111011" => data <= "000000";
				when "001110101000111100" => data <= "000000";
				when "001110101000111101" => data <= "000000";
				when "001110101000111110" => data <= "000000";
				when "001110101000111111" => data <= "000000";
				when "001110101001000000" => data <= "000000";
				when "001110101001000001" => data <= "000000";
				when "001110101001000010" => data <= "000000";
				when "001110101001000011" => data <= "000000";
				when "001110101001000100" => data <= "000000";
				when "001110101001000101" => data <= "000000";
				when "001110101001000110" => data <= "000000";
				when "001110101001000111" => data <= "000000";
				when "001110101001001000" => data <= "000000";
				when "001110101001001001" => data <= "000000";
				when "001110101001001010" => data <= "000000";
				when "001110101001001011" => data <= "000000";
				when "001110101001001100" => data <= "000000";
				when "001110101001001101" => data <= "000000";
				when "001110101001001110" => data <= "000000";
				when "001110101001001111" => data <= "000000";
				when "001110101001010000" => data <= "000000";
				when "001110101001010001" => data <= "000000";
				when "001110101001010010" => data <= "000000";
				when "001110101001010011" => data <= "000000";
				when "001110101001010100" => data <= "000000";
				when "001110101001010101" => data <= "000000";
				when "001110101001010110" => data <= "000000";
				when "001110101001010111" => data <= "000000";
				when "001110101001011000" => data <= "000000";
				when "001110101001011001" => data <= "000000";
				when "001110101001011010" => data <= "000000";
				when "001110101001011011" => data <= "000000";
				when "001110101001011100" => data <= "000000";
				when "001110101001011101" => data <= "000000";
				when "001110101001011110" => data <= "000000";
				when "001110101001011111" => data <= "000000";
				when "001110101001100000" => data <= "000000";
				when "001110101001100001" => data <= "000000";
				when "001110101001100010" => data <= "000000";
				when "001110101001100011" => data <= "000000";
				when "001110101001100100" => data <= "000000";
				when "001110101001100101" => data <= "000000";
				when "001110101001100110" => data <= "000000";
				when "001110101001100111" => data <= "000000";
				when "001110101001101000" => data <= "000000";
				when "001110101001101001" => data <= "000000";
				when "001110101001101010" => data <= "000000";
				when "001110101001101011" => data <= "000000";
				when "001110101001101100" => data <= "000000";
				when "001110101001101101" => data <= "000000";
				when "001110101001101110" => data <= "000000";
				when "001110101001101111" => data <= "000000";
				when "001110101001110000" => data <= "000000";
				when "001110101001110001" => data <= "000000";
				when "001110101001110010" => data <= "000000";
				when "001110101001110011" => data <= "000000";
				when "001110101001110100" => data <= "000000";
				when "001110101001110101" => data <= "000000";
				when "001110101001110110" => data <= "000000";
				when "001110101001110111" => data <= "000000";
				when "001110101001111000" => data <= "000000";
				when "001110101001111001" => data <= "000000";
				when "001110101001111010" => data <= "000000";
				when "001110101001111011" => data <= "000000";
				when "001110101001111100" => data <= "000000";
				when "001110101001111101" => data <= "000000";
				when "001110101001111110" => data <= "000000";
				when "001110101001111111" => data <= "000000";
				when "001110101010000000" => data <= "000000";
				when "001110101010000001" => data <= "000000";
				when "001110101010000010" => data <= "000000";
				when "001110101010000011" => data <= "000000";
				when "001110101010000100" => data <= "000000";
				when "001110101010000101" => data <= "000000";
				when "001110101010000110" => data <= "000000";
				when "001110101010000111" => data <= "000000";
				when "001110101010001000" => data <= "000000";
				when "001110101010001001" => data <= "000000";
				when "001110101010001010" => data <= "000000";
				when "001110101010001011" => data <= "000000";
				when "001110101010001100" => data <= "000000";
				when "001110101010001101" => data <= "000000";
				when "001110101010001110" => data <= "000000";
				when "001110101010001111" => data <= "000000";
				when "001110101010010000" => data <= "000000";
				when "001110101010010001" => data <= "000000";
				when "001110101010010010" => data <= "000000";
				when "001110101010010011" => data <= "000000";
				when "001110101010010100" => data <= "000000";
				when "001110101010010101" => data <= "000000";
				when "001110101010010110" => data <= "000000";
				when "001110101010010111" => data <= "000000";
				when "001110101010011000" => data <= "000000";
				when "001110101010011001" => data <= "000000";
				when "001110101010011010" => data <= "000000";
				when "001110101010011011" => data <= "000000";
				when "001110101010011100" => data <= "000000";
				when "001110101010011101" => data <= "000000";
				when "001110101010011110" => data <= "000000";
				when "001110101010011111" => data <= "000000";
				when "001110110000000000" => data <= "000000";
				when "001110110000000001" => data <= "000000";
				when "001110110000000010" => data <= "000000";
				when "001110110000000011" => data <= "000000";
				when "001110110000000100" => data <= "000000";
				when "001110110000000101" => data <= "000000";
				when "001110110000000110" => data <= "000000";
				when "001110110000000111" => data <= "000000";
				when "001110110000001000" => data <= "000000";
				when "001110110000001001" => data <= "000000";
				when "001110110000001010" => data <= "000000";
				when "001110110000001011" => data <= "000000";
				when "001110110000001100" => data <= "000000";
				when "001110110000001101" => data <= "000000";
				when "001110110000001110" => data <= "000000";
				when "001110110000001111" => data <= "000000";
				when "001110110000010000" => data <= "000000";
				when "001110110000010001" => data <= "000000";
				when "001110110000010010" => data <= "000000";
				when "001110110000010011" => data <= "000000";
				when "001110110000010100" => data <= "000000";
				when "001110110000010101" => data <= "000000";
				when "001110110000010110" => data <= "000000";
				when "001110110000010111" => data <= "000000";
				when "001110110000011000" => data <= "000000";
				when "001110110000011001" => data <= "000000";
				when "001110110000011010" => data <= "000000";
				when "001110110000011011" => data <= "000000";
				when "001110110000011100" => data <= "000000";
				when "001110110000011101" => data <= "000000";
				when "001110110000011110" => data <= "000000";
				when "001110110000011111" => data <= "000000";
				when "001110110000100000" => data <= "000000";
				when "001110110000100001" => data <= "000000";
				when "001110110000100010" => data <= "000000";
				when "001110110000100011" => data <= "000000";
				when "001110110000100100" => data <= "000000";
				when "001110110000100101" => data <= "000000";
				when "001110110000100110" => data <= "000000";
				when "001110110000100111" => data <= "000000";
				when "001110110000101000" => data <= "000000";
				when "001110110000101001" => data <= "000000";
				when "001110110000101010" => data <= "000000";
				when "001110110000101011" => data <= "000000";
				when "001110110000101100" => data <= "000000";
				when "001110110000101101" => data <= "000000";
				when "001110110000101110" => data <= "000000";
				when "001110110000101111" => data <= "000000";
				when "001110110000110000" => data <= "000000";
				when "001110110000110001" => data <= "000000";
				when "001110110000110010" => data <= "000000";
				when "001110110000110011" => data <= "000000";
				when "001110110000110100" => data <= "000000";
				when "001110110000110101" => data <= "000000";
				when "001110110000110110" => data <= "000000";
				when "001110110000110111" => data <= "000000";
				when "001110110000111000" => data <= "000000";
				when "001110110000111001" => data <= "000000";
				when "001110110000111010" => data <= "000000";
				when "001110110000111011" => data <= "000000";
				when "001110110000111100" => data <= "000000";
				when "001110110000111101" => data <= "000000";
				when "001110110000111110" => data <= "000000";
				when "001110110000111111" => data <= "000000";
				when "001110110001000000" => data <= "000000";
				when "001110110001000001" => data <= "000000";
				when "001110110001000010" => data <= "000000";
				when "001110110001000011" => data <= "000000";
				when "001110110001000100" => data <= "000000";
				when "001110110001000101" => data <= "000000";
				when "001110110001000110" => data <= "000000";
				when "001110110001000111" => data <= "000000";
				when "001110110001001000" => data <= "000000";
				when "001110110001001001" => data <= "000000";
				when "001110110001001010" => data <= "000000";
				when "001110110001001011" => data <= "000000";
				when "001110110001001100" => data <= "000000";
				when "001110110001001101" => data <= "000000";
				when "001110110001001110" => data <= "000000";
				when "001110110001001111" => data <= "000000";
				when "001110110001010000" => data <= "000000";
				when "001110110001010001" => data <= "000000";
				when "001110110001010010" => data <= "000000";
				when "001110110001010011" => data <= "000000";
				when "001110110001010100" => data <= "000000";
				when "001110110001010101" => data <= "000000";
				when "001110110001010110" => data <= "000000";
				when "001110110001010111" => data <= "000000";
				when "001110110001011000" => data <= "000000";
				when "001110110001011001" => data <= "000000";
				when "001110110001011010" => data <= "000000";
				when "001110110001011011" => data <= "000000";
				when "001110110001011100" => data <= "000000";
				when "001110110001011101" => data <= "000000";
				when "001110110001011110" => data <= "000000";
				when "001110110001011111" => data <= "000000";
				when "001110110001100000" => data <= "000000";
				when "001110110001100001" => data <= "000000";
				when "001110110001100010" => data <= "000000";
				when "001110110001100011" => data <= "000000";
				when "001110110001100100" => data <= "000000";
				when "001110110001100101" => data <= "000000";
				when "001110110001100110" => data <= "000000";
				when "001110110001100111" => data <= "000000";
				when "001110110001101000" => data <= "000000";
				when "001110110001101001" => data <= "000000";
				when "001110110001101010" => data <= "000000";
				when "001110110001101011" => data <= "000000";
				when "001110110001101100" => data <= "000000";
				when "001110110001101101" => data <= "000000";
				when "001110110001101110" => data <= "000000";
				when "001110110001101111" => data <= "000000";
				when "001110110001110000" => data <= "000000";
				when "001110110001110001" => data <= "000000";
				when "001110110001110010" => data <= "000000";
				when "001110110001110011" => data <= "000000";
				when "001110110001110100" => data <= "000000";
				when "001110110001110101" => data <= "000000";
				when "001110110001110110" => data <= "000000";
				when "001110110001110111" => data <= "000000";
				when "001110110001111000" => data <= "000000";
				when "001110110001111001" => data <= "000000";
				when "001110110001111010" => data <= "000000";
				when "001110110001111011" => data <= "000000";
				when "001110110001111100" => data <= "000000";
				when "001110110001111101" => data <= "000000";
				when "001110110001111110" => data <= "000000";
				when "001110110001111111" => data <= "000000";
				when "001110110010000000" => data <= "000000";
				when "001110110010000001" => data <= "000000";
				when "001110110010000010" => data <= "000000";
				when "001110110010000011" => data <= "000000";
				when "001110110010000100" => data <= "000000";
				when "001110110010000101" => data <= "000000";
				when "001110110010000110" => data <= "000000";
				when "001110110010000111" => data <= "000000";
				when "001110110010001000" => data <= "000000";
				when "001110110010001001" => data <= "000000";
				when "001110110010001010" => data <= "000000";
				when "001110110010001011" => data <= "000000";
				when "001110110010001100" => data <= "000000";
				when "001110110010001101" => data <= "000000";
				when "001110110010001110" => data <= "000000";
				when "001110110010001111" => data <= "000000";
				when "001110110010010000" => data <= "000000";
				when "001110110010010001" => data <= "000000";
				when "001110110010010010" => data <= "000000";
				when "001110110010010011" => data <= "000000";
				when "001110110010010100" => data <= "000000";
				when "001110110010010101" => data <= "000000";
				when "001110110010010110" => data <= "000000";
				when "001110110010010111" => data <= "000000";
				when "001110110010011000" => data <= "000000";
				when "001110110010011001" => data <= "000000";
				when "001110110010011010" => data <= "000000";
				when "001110110010011011" => data <= "000000";
				when "001110110010011100" => data <= "000000";
				when "001110110010011101" => data <= "000000";
				when "001110110010011110" => data <= "000000";
				when "001110110010011111" => data <= "000000";
				when "001110111000000000" => data <= "000000";
				when "001110111000000001" => data <= "000000";
				when "001110111000000010" => data <= "000000";
				when "001110111000000011" => data <= "000000";
				when "001110111000000100" => data <= "000000";
				when "001110111000000101" => data <= "000000";
				when "001110111000000110" => data <= "000000";
				when "001110111000000111" => data <= "000000";
				when "001110111000001000" => data <= "000000";
				when "001110111000001001" => data <= "000000";
				when "001110111000001010" => data <= "000000";
				when "001110111000001011" => data <= "000000";
				when "001110111000001100" => data <= "000000";
				when "001110111000001101" => data <= "000000";
				when "001110111000001110" => data <= "000000";
				when "001110111000001111" => data <= "000000";
				when "001110111000010000" => data <= "000000";
				when "001110111000010001" => data <= "000000";
				when "001110111000010010" => data <= "000000";
				when "001110111000010011" => data <= "000000";
				when "001110111000010100" => data <= "000000";
				when "001110111000010101" => data <= "000000";
				when "001110111000010110" => data <= "000000";
				when "001110111000010111" => data <= "000000";
				when "001110111000011000" => data <= "000000";
				when "001110111000011001" => data <= "000000";
				when "001110111000011010" => data <= "000000";
				when "001110111000011011" => data <= "000000";
				when "001110111000011100" => data <= "000000";
				when "001110111000011101" => data <= "000000";
				when "001110111000011110" => data <= "000000";
				when "001110111000011111" => data <= "000000";
				when "001110111000100000" => data <= "000000";
				when "001110111000100001" => data <= "000000";
				when "001110111000100010" => data <= "000000";
				when "001110111000100011" => data <= "000000";
				when "001110111000100100" => data <= "000000";
				when "001110111000100101" => data <= "000000";
				when "001110111000100110" => data <= "000000";
				when "001110111000100111" => data <= "000000";
				when "001110111000101000" => data <= "000000";
				when "001110111000101001" => data <= "000000";
				when "001110111000101010" => data <= "000000";
				when "001110111000101011" => data <= "000000";
				when "001110111000101100" => data <= "000000";
				when "001110111000101101" => data <= "000000";
				when "001110111000101110" => data <= "000000";
				when "001110111000101111" => data <= "000000";
				when "001110111000110000" => data <= "000000";
				when "001110111000110001" => data <= "000000";
				when "001110111000110010" => data <= "000000";
				when "001110111000110011" => data <= "000000";
				when "001110111000110100" => data <= "000000";
				when "001110111000110101" => data <= "000000";
				when "001110111000110110" => data <= "000000";
				when "001110111000110111" => data <= "000000";
				when "001110111000111000" => data <= "000000";
				when "001110111000111001" => data <= "000000";
				when "001110111000111010" => data <= "000000";
				when "001110111000111011" => data <= "000000";
				when "001110111000111100" => data <= "000000";
				when "001110111000111101" => data <= "000000";
				when "001110111000111110" => data <= "000000";
				when "001110111000111111" => data <= "000000";
				when "001110111001000000" => data <= "000000";
				when "001110111001000001" => data <= "000000";
				when "001110111001000010" => data <= "000000";
				when "001110111001000011" => data <= "000000";
				when "001110111001000100" => data <= "000000";
				when "001110111001000101" => data <= "000000";
				when "001110111001000110" => data <= "000000";
				when "001110111001000111" => data <= "000000";
				when "001110111001001000" => data <= "000000";
				when "001110111001001001" => data <= "000000";
				when "001110111001001010" => data <= "000000";
				when "001110111001001011" => data <= "000000";
				when "001110111001001100" => data <= "000000";
				when "001110111001001101" => data <= "000000";
				when "001110111001001110" => data <= "000000";
				when "001110111001001111" => data <= "000000";
				when "001110111001010000" => data <= "000000";
				when "001110111001010001" => data <= "000000";
				when "001110111001010010" => data <= "000000";
				when "001110111001010011" => data <= "000000";
				when "001110111001010100" => data <= "000000";
				when "001110111001010101" => data <= "000000";
				when "001110111001010110" => data <= "000000";
				when "001110111001010111" => data <= "000000";
				when "001110111001011000" => data <= "000000";
				when "001110111001011001" => data <= "000000";
				when "001110111001011010" => data <= "000000";
				when "001110111001011011" => data <= "000000";
				when "001110111001011100" => data <= "000000";
				when "001110111001011101" => data <= "000000";
				when "001110111001011110" => data <= "000000";
				when "001110111001011111" => data <= "000000";
				when "001110111001100000" => data <= "000000";
				when "001110111001100001" => data <= "000000";
				when "001110111001100010" => data <= "000000";
				when "001110111001100011" => data <= "000000";
				when "001110111001100100" => data <= "000000";
				when "001110111001100101" => data <= "000000";
				when "001110111001100110" => data <= "000000";
				when "001110111001100111" => data <= "000000";
				when "001110111001101000" => data <= "000000";
				when "001110111001101001" => data <= "000000";
				when "001110111001101010" => data <= "000000";
				when "001110111001101011" => data <= "000000";
				when "001110111001101100" => data <= "000000";
				when "001110111001101101" => data <= "000000";
				when "001110111001101110" => data <= "000000";
				when "001110111001101111" => data <= "000000";
				when "001110111001110000" => data <= "000000";
				when "001110111001110001" => data <= "000000";
				when "001110111001110010" => data <= "000000";
				when "001110111001110011" => data <= "000000";
				when "001110111001110100" => data <= "000000";
				when "001110111001110101" => data <= "000000";
				when "001110111001110110" => data <= "000000";
				when "001110111001110111" => data <= "000000";
				when "001110111001111000" => data <= "000000";
				when "001110111001111001" => data <= "000000";
				when "001110111001111010" => data <= "000000";
				when "001110111001111011" => data <= "000000";
				when "001110111001111100" => data <= "000000";
				when "001110111001111101" => data <= "000000";
				when "001110111001111110" => data <= "000000";
				when "001110111001111111" => data <= "000000";
				when "001110111010000000" => data <= "000000";
				when "001110111010000001" => data <= "000000";
				when "001110111010000010" => data <= "000000";
				when "001110111010000011" => data <= "000000";
				when "001110111010000100" => data <= "000000";
				when "001110111010000101" => data <= "000000";
				when "001110111010000110" => data <= "000000";
				when "001110111010000111" => data <= "000000";
				when "001110111010001000" => data <= "000000";
				when "001110111010001001" => data <= "000000";
				when "001110111010001010" => data <= "000000";
				when "001110111010001011" => data <= "000000";
				when "001110111010001100" => data <= "000000";
				when "001110111010001101" => data <= "000000";
				when "001110111010001110" => data <= "000000";
				when "001110111010001111" => data <= "000000";
				when "001110111010010000" => data <= "000000";
				when "001110111010010001" => data <= "000000";
				when "001110111010010010" => data <= "000000";
				when "001110111010010011" => data <= "000000";
				when "001110111010010100" => data <= "000000";
				when "001110111010010101" => data <= "000000";
				when "001110111010010110" => data <= "000000";
				when "001110111010010111" => data <= "000000";
				when "001110111010011000" => data <= "000000";
				when "001110111010011001" => data <= "000000";
				when "001110111010011010" => data <= "000000";
				when "001110111010011011" => data <= "000000";
				when "001110111010011100" => data <= "000000";
				when "001110111010011101" => data <= "000000";
				when "001110111010011110" => data <= "000000";
				when "001110111010011111" => data <= "000000";
				when others => data <= "000000";
			end case;
              		end if; 
              	end process; 
              end;