library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity score_disp is 
 	port(
		outglobal_o : in std_logic;
		addr_x : in std_logic_vector(7 downto 0);
		addr_y : in std_logic_vector(7 downto 0);
		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
	);
end;

architecture sim of score_disp is
signal addr : std_logic_vector(15 downto 0);

begin
	addr (15 downto 8) <= addr_x;
	addr (7 downto 0) <= addr_y;
	process(outglobal_o) begin
		if rising_edge(outglobal_o) then
			case addr is
				when "0000000000000000" => data <= "000001";
				when "0000000000000001" => data <= "111111";
				when "0000000000000010" => data <= "111111";
				when "0000000000000011" => data <= "111111";
				when "0000000000000100" => data <= "111111";
				when "0000000000000101" => data <= "000001";
				when "0000000000000110" => data <= "111111";
				when "0000000000000111" => data <= "111111";
				when "0000000000001000" => data <= "111111";
				when "0000000000001001" => data <= "111111";
				when "0000000000001010" => data <= "000001";
				when "0000000000001011" => data <= "111111";
				when "0000000000001100" => data <= "111111";
				when "0000000000001101" => data <= "111111";
				when "0000000000001110" => data <= "111111";
				when "0000000000001111" => data <= "111111";
				when "0000000000010000" => data <= "000001";
				when "0000000000010001" => data <= "111111";
				when "0000000000010010" => data <= "111111";
				when "0000000000010011" => data <= "111111";
				when "0000000000010100" => data <= "111111";
				when "0000000000010101" => data <= "000001";
				when "0000000000010110" => data <= "000001";
				when "0000000000010111" => data <= "111111";
				when "0000000000011000" => data <= "111111";
				when "0000000000011001" => data <= "111111";
				when "0000000000011010" => data <= "111111";
				when "0000000000011011" => data <= "000001";
				when "0000000000011100" => data <= "000001";
				when "0000000000011101" => data <= "000001";
				when "0000000100000000" => data <= "000001";
				when "0000000100000001" => data <= "111111";
				when "0000000100000010" => data <= "000001";
				when "0000000100000011" => data <= "000001";
				when "0000000100000100" => data <= "000001";
				when "0000000100000101" => data <= "000001";
				when "0000000100000110" => data <= "111111";
				when "0000000100000111" => data <= "000001";
				when "0000000100001000" => data <= "000001";
				when "0000000100001001" => data <= "000001";
				when "0000000100001010" => data <= "000001";
				when "0000000100001011" => data <= "111111";
				when "0000000100001100" => data <= "000001";
				when "0000000100001101" => data <= "000001";
				when "0000000100001110" => data <= "000001";
				when "0000000100001111" => data <= "111111";
				when "0000000100010000" => data <= "000001";
				when "0000000100010001" => data <= "111111";
				when "0000000100010010" => data <= "000001";
				when "0000000100010011" => data <= "000001";
				when "0000000100010100" => data <= "000001";
				when "0000000100010101" => data <= "111111";
				when "0000000100010110" => data <= "000001";
				when "0000000100010111" => data <= "111111";
				when "0000000100011000" => data <= "000001";
				when "0000000100011001" => data <= "000001";
				when "0000000100011010" => data <= "000001";
				when "0000000100011011" => data <= "000001";
				when "0000000100011100" => data <= "000001";
				when "0000000100011101" => data <= "000001";
				when "0000001000000000" => data <= "000001";
				when "0000001000000001" => data <= "111111";
				when "0000001000000010" => data <= "000001";
				when "0000001000000011" => data <= "000001";
				when "0000001000000100" => data <= "000001";
				when "0000001000000101" => data <= "000001";
				when "0000001000000110" => data <= "111111";
				when "0000001000000111" => data <= "000001";
				when "0000001000001000" => data <= "000001";
				when "0000001000001001" => data <= "000001";
				when "0000001000001010" => data <= "000001";
				when "0000001000001011" => data <= "111111";
				when "0000001000001100" => data <= "000001";
				when "0000001000001101" => data <= "000001";
				when "0000001000001110" => data <= "000001";
				when "0000001000001111" => data <= "111111";
				when "0000001000010000" => data <= "000001";
				when "0000001000010001" => data <= "111111";
				when "0000001000010010" => data <= "000001";
				when "0000001000010011" => data <= "000001";
				when "0000001000010100" => data <= "000001";
				when "0000001000010101" => data <= "111111";
				when "0000001000010110" => data <= "000001";
				when "0000001000010111" => data <= "111111";
				when "0000001000011000" => data <= "000001";
				when "0000001000011001" => data <= "000001";
				when "0000001000011010" => data <= "000001";
				when "0000001000011011" => data <= "000001";
				when "0000001000011100" => data <= "111111";
				when "0000001000011101" => data <= "000001";
				when "0000001100000000" => data <= "000001";
				when "0000001100000001" => data <= "111111";
				when "0000001100000010" => data <= "111111";
				when "0000001100000011" => data <= "111111";
				when "0000001100000100" => data <= "111111";
				when "0000001100000101" => data <= "000001";
				when "0000001100000110" => data <= "111111";
				when "0000001100000111" => data <= "000001";
				when "0000001100001000" => data <= "000001";
				when "0000001100001001" => data <= "000001";
				when "0000001100001010" => data <= "000001";
				when "0000001100001011" => data <= "111111";
				when "0000001100001100" => data <= "000001";
				when "0000001100001101" => data <= "000001";
				when "0000001100001110" => data <= "000001";
				when "0000001100001111" => data <= "111111";
				when "0000001100010000" => data <= "000001";
				when "0000001100010001" => data <= "111111";
				when "0000001100010010" => data <= "000001";
				when "0000001100010011" => data <= "000001";
				when "0000001100010100" => data <= "000001";
				when "0000001100010101" => data <= "111111";
				when "0000001100010110" => data <= "000001";
				when "0000001100010111" => data <= "111111";
				when "0000001100011000" => data <= "111111";
				when "0000001100011001" => data <= "111111";
				when "0000001100011010" => data <= "000001";
				when "0000001100011011" => data <= "000001";
				when "0000001100011100" => data <= "000001";
				when "0000001100011101" => data <= "000001";
				when "0000010000000000" => data <= "000001";
				when "0000010000000001" => data <= "000001";
				when "0000010000000010" => data <= "000001";
				when "0000010000000011" => data <= "000001";
				when "0000010000000100" => data <= "111111";
				when "0000010000000101" => data <= "000001";
				when "0000010000000110" => data <= "111111";
				when "0000010000000111" => data <= "000001";
				when "0000010000001000" => data <= "000001";
				when "0000010000001001" => data <= "000001";
				when "0000010000001010" => data <= "000001";
				when "0000010000001011" => data <= "111111";
				when "0000010000001100" => data <= "000001";
				when "0000010000001101" => data <= "000001";
				when "0000010000001110" => data <= "000001";
				when "0000010000001111" => data <= "111111";
				when "0000010000010000" => data <= "000001";
				when "0000010000010001" => data <= "111111";
				when "0000010000010010" => data <= "111111";
				when "0000010000010011" => data <= "111111";
				when "0000010000010100" => data <= "111111";
				when "0000010000010101" => data <= "000001";
				when "0000010000010110" => data <= "000001";
				when "0000010000010111" => data <= "111111";
				when "0000010000011000" => data <= "000001";
				when "0000010000011001" => data <= "000001";
				when "0000010000011010" => data <= "000001";
				when "0000010000011011" => data <= "000001";
				when "0000010000011100" => data <= "000001";
				when "0000010000011101" => data <= "000001";
				when "0000010100000000" => data <= "000001";
				when "0000010100000001" => data <= "000001";
				when "0000010100000010" => data <= "000001";
				when "0000010100000011" => data <= "000001";
				when "0000010100000100" => data <= "111111";
				when "0000010100000101" => data <= "000001";
				when "0000010100000110" => data <= "111111";
				when "0000010100000111" => data <= "000001";
				when "0000010100001000" => data <= "000001";
				when "0000010100001001" => data <= "000001";
				when "0000010100001010" => data <= "000001";
				when "0000010100001011" => data <= "111111";
				when "0000010100001100" => data <= "000001";
				when "0000010100001101" => data <= "000001";
				when "0000010100001110" => data <= "000001";
				when "0000010100001111" => data <= "111111";
				when "0000010100010000" => data <= "000001";
				when "0000010100010001" => data <= "111111";
				when "0000010100010010" => data <= "000001";
				when "0000010100010011" => data <= "000001";
				when "0000010100010100" => data <= "000001";
				when "0000010100010101" => data <= "111111";
				when "0000010100010110" => data <= "000001";
				when "0000010100010111" => data <= "111111";
				when "0000010100011000" => data <= "000001";
				when "0000010100011001" => data <= "000001";
				when "0000010100011010" => data <= "000001";
				when "0000010100011011" => data <= "000001";
				when "0000010100011100" => data <= "111111";
				when "0000010100011101" => data <= "000001";
				when "0000011000000000" => data <= "000001";
				when "0000011000000001" => data <= "000001";
				when "0000011000000010" => data <= "000001";
				when "0000011000000011" => data <= "000001";
				when "0000011000000100" => data <= "111111";
				when "0000011000000101" => data <= "000001";
				when "0000011000000110" => data <= "111111";
				when "0000011000000111" => data <= "000001";
				when "0000011000001000" => data <= "000001";
				when "0000011000001001" => data <= "000001";
				when "0000011000001010" => data <= "000001";
				when "0000011000001011" => data <= "111111";
				when "0000011000001100" => data <= "000001";
				when "0000011000001101" => data <= "000001";
				when "0000011000001110" => data <= "000001";
				when "0000011000001111" => data <= "111111";
				when "0000011000010000" => data <= "000001";
				when "0000011000010001" => data <= "111111";
				when "0000011000010010" => data <= "000001";
				when "0000011000010011" => data <= "000001";
				when "0000011000010100" => data <= "000001";
				when "0000011000010101" => data <= "111111";
				when "0000011000010110" => data <= "000001";
				when "0000011000010111" => data <= "111111";
				when "0000011000011000" => data <= "000001";
				when "0000011000011001" => data <= "000001";
				when "0000011000011010" => data <= "000001";
				when "0000011000011011" => data <= "000001";
				when "0000011000011100" => data <= "000001";
				when "0000011000011101" => data <= "000001";
				when "0000011100000000" => data <= "000001";
				when "0000011100000001" => data <= "111111";
				when "0000011100000010" => data <= "111111";
				when "0000011100000011" => data <= "111111";
				when "0000011100000100" => data <= "111111";
				when "0000011100000101" => data <= "000001";
				when "0000011100000110" => data <= "111111";
				when "0000011100000111" => data <= "111111";
				when "0000011100001000" => data <= "111111";
				when "0000011100001001" => data <= "111111";
				when "0000011100001010" => data <= "000001";
				when "0000011100001011" => data <= "111111";
				when "0000011100001100" => data <= "111111";
				when "0000011100001101" => data <= "111111";
				when "0000011100001110" => data <= "111111";
				when "0000011100001111" => data <= "111111";
				when "0000011100010000" => data <= "000001";
				when "0000011100010001" => data <= "111111";
				when "0000011100010010" => data <= "000001";
				when "0000011100010011" => data <= "000001";
				when "0000011100010100" => data <= "000001";
				when "0000011100010101" => data <= "111111";
				when "0000011100010110" => data <= "000001";
				when "0000011100010111" => data <= "111111";
				when "0000011100011000" => data <= "111111";
				when "0000011100011001" => data <= "111111";
				when "0000011100011010" => data <= "111111";
				when "0000011100011011" => data <= "000001";
				when "0000011100011100" => data <= "000001";
				when "0000011100011101" => data <= "000001";
				when others => data <= "010001";
			end case;
		end if; 
	end process; 
end;