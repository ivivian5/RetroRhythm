library IEEE;
                use IEEE.std_logic_1164.all;
                use IEEE.numeric_std.all;

entity endscreen is 
                 	port(
                		outglobal_o : in std_logic;
                		addr_x : in std_logic_vector(7 downto 0);
                		addr_y : in std_logic_vector(7 downto 0);
                		data : out std_logic_vector(5 downto 0) -- 6-bit words, RRGGBB
                	);
                end;

                architecture sim of endscreen is
                signal addr : std_logic_vector(15 downto 0);

                begin
                	addr (15 downto 8) <= addr_x;
                	addr (7 downto 0) <= addr_y;
                	process(outglobal_o) begin
                		if rising_edge(outglobal_o) then
                			case addr is
				when "0001100100101001" => data <= "111111";
				when "0001100100101010" => data <= "111111";
				when "0001100100101011" => data <= "111111";
				when "0001100100101100" => data <= "111111";
				when "0001100100101101" => data <= "111111";
				when "0001100100101110" => data <= "111111";
				when "0001100100101111" => data <= "111111";
				when "0001100100110000" => data <= "111111";
				when "0001100100110001" => data <= "111111";
				when "0001100100110010" => data <= "111111";
				when "0001100100110011" => data <= "111111";
				when "0001100100111100" => data <= "111111";
				when "0001100100111101" => data <= "111111";
				when "0001100100111110" => data <= "111111";
				when "0001100100111111" => data <= "111111";
				when "0001100101000000" => data <= "111111";
				when "0001100101000001" => data <= "111111";
				when "0001100101000010" => data <= "111111";
				when "0001100101000011" => data <= "111111";
				when "0001100101000100" => data <= "111111";
				when "0001100101000101" => data <= "111111";
				when "0001100101000110" => data <= "111111";
				when "0001100101010000" => data <= "111111";
				when "0001100101010001" => data <= "111111";
				when "0001100101010010" => data <= "111111";
				when "0001100101010011" => data <= "111111";
				when "0001100101011100" => data <= "111111";
				when "0001100101011101" => data <= "111111";
				when "0001100101011110" => data <= "111111";
				when "0001100101011111" => data <= "111111";
				when "0001100101101001" => data <= "111111";
				when "0001100101101010" => data <= "111111";
				when "0001100101101011" => data <= "111111";
				when "0001100101101100" => data <= "111111";
				when "0001100101101101" => data <= "111111";
				when "0001100101101110" => data <= "111111";
				when "0001100101101111" => data <= "111111";
				when "0001100101110000" => data <= "111111";
				when "0001100101110001" => data <= "111111";
				when "0001100101110010" => data <= "111111";
				when "0001100101110011" => data <= "111111";
				when "0001101000101000" => data <= "111111";
				when "0001101000101001" => data <= "100110";
				when "0001101000101010" => data <= "010110";
				when "0001101000101011" => data <= "010110";
				when "0001101000101100" => data <= "100110";
				when "0001101000101101" => data <= "010110";
				when "0001101000101110" => data <= "010110";
				when "0001101000101111" => data <= "010110";
				when "0001101000110000" => data <= "010110";
				when "0001101000110001" => data <= "010110";
				when "0001101000110010" => data <= "010110";
				when "0001101000110011" => data <= "111111";
				when "0001101000111011" => data <= "111111";
				when "0001101000111100" => data <= "100110";
				when "0001101000111101" => data <= "100110";
				when "0001101000111110" => data <= "100110";
				when "0001101000111111" => data <= "100110";
				when "0001101001000000" => data <= "100110";
				when "0001101001000001" => data <= "010110";
				when "0001101001000010" => data <= "100110";
				when "0001101001000011" => data <= "100110";
				when "0001101001000100" => data <= "100110";
				when "0001101001000101" => data <= "100110";
				when "0001101001000110" => data <= "100110";
				when "0001101001000111" => data <= "111111";
				when "0001101001001111" => data <= "111111";
				when "0001101001010000" => data <= "010110";
				when "0001101001010001" => data <= "100110";
				when "0001101001010010" => data <= "100110";
				when "0001101001010011" => data <= "100110";
				when "0001101001010100" => data <= "111111";
				when "0001101001011011" => data <= "111111";
				when "0001101001011100" => data <= "100110";
				when "0001101001011101" => data <= "100110";
				when "0001101001011110" => data <= "100110";
				when "0001101001011111" => data <= "100110";
				when "0001101001100000" => data <= "111111";
				when "0001101001101000" => data <= "111111";
				when "0001101001101001" => data <= "100110";
				when "0001101001101010" => data <= "100110";
				when "0001101001101011" => data <= "100110";
				when "0001101001101100" => data <= "100110";
				when "0001101001101101" => data <= "100110";
				when "0001101001101110" => data <= "100110";
				when "0001101001101111" => data <= "100110";
				when "0001101001110000" => data <= "100110";
				when "0001101001110001" => data <= "100110";
				when "0001101001110010" => data <= "100110";
				when "0001101001110011" => data <= "100110";
				when "0001101001110100" => data <= "111111";
				when "0001101100101000" => data <= "111111";
				when "0001101100101001" => data <= "100110";
				when "0001101100101010" => data <= "100110";
				when "0001101100101011" => data <= "100110";
				when "0001101100101100" => data <= "111111";
				when "0001101100101101" => data <= "111111";
				when "0001101100101110" => data <= "111111";
				when "0001101100101111" => data <= "111111";
				when "0001101100110000" => data <= "111111";
				when "0001101100110001" => data <= "111111";
				when "0001101100110010" => data <= "111111";
				when "0001101100110011" => data <= "111111";
				when "0001101100111011" => data <= "111111";
				when "0001101100111100" => data <= "100110";
				when "0001101100111101" => data <= "100111";
				when "0001101100111110" => data <= "100110";
				when "0001101100111111" => data <= "100110";
				when "0001101101000000" => data <= "100110";
				when "0001101101000001" => data <= "100110";
				when "0001101101000010" => data <= "100110";
				when "0001101101000011" => data <= "100110";
				when "0001101101000100" => data <= "100110";
				when "0001101101000101" => data <= "100110";
				when "0001101101000110" => data <= "100110";
				when "0001101101000111" => data <= "111111";
				when "0001101101001111" => data <= "111111";
				when "0001101101010000" => data <= "100110";
				when "0001101101010001" => data <= "100111";
				when "0001101101010010" => data <= "100111";
				when "0001101101010011" => data <= "100111";
				when "0001101101010100" => data <= "100110";
				when "0001101101010101" => data <= "111111";
				when "0001101101011010" => data <= "111111";
				when "0001101101011011" => data <= "100110";
				when "0001101101011100" => data <= "100110";
				when "0001101101011101" => data <= "100110";
				when "0001101101011110" => data <= "100110";
				when "0001101101011111" => data <= "100110";
				when "0001101101100000" => data <= "111111";
				when "0001101101101000" => data <= "111111";
				when "0001101101101001" => data <= "100110";
				when "0001101101101010" => data <= "100110";
				when "0001101101101011" => data <= "100110";
				when "0001101101101100" => data <= "100110";
				when "0001101101101101" => data <= "100110";
				when "0001101101101110" => data <= "100110";
				when "0001101101101111" => data <= "010110";
				when "0001101101110000" => data <= "100110";
				when "0001101101110001" => data <= "100110";
				when "0001101101110010" => data <= "010110";
				when "0001101101110011" => data <= "010110";
				when "0001101101110100" => data <= "111111";
				when "0001110000101000" => data <= "111111";
				when "0001110000101001" => data <= "100110";
				when "0001110000101010" => data <= "100110";
				when "0001110000101011" => data <= "100110";
				when "0001110000101100" => data <= "111111";
				when "0001110000111011" => data <= "111111";
				when "0001110000111100" => data <= "100110";
				when "0001110000111101" => data <= "100111";
				when "0001110000111110" => data <= "100110";
				when "0001110000111111" => data <= "100110";
				when "0001110001000000" => data <= "100110";
				when "0001110001000001" => data <= "100110";
				when "0001110001000010" => data <= "100110";
				when "0001110001000011" => data <= "100110";
				when "0001110001000100" => data <= "100110";
				when "0001110001000101" => data <= "100110";
				when "0001110001000110" => data <= "100110";
				when "0001110001000111" => data <= "111111";
				when "0001110001001111" => data <= "111111";
				when "0001110001010000" => data <= "100110";
				when "0001110001010001" => data <= "100111";
				when "0001110001010010" => data <= "100111";
				when "0001110001010011" => data <= "100111";
				when "0001110001010100" => data <= "100110";
				when "0001110001010101" => data <= "111111";
				when "0001110001011010" => data <= "111111";
				when "0001110001011011" => data <= "100110";
				when "0001110001011100" => data <= "100110";
				when "0001110001011101" => data <= "100110";
				when "0001110001011110" => data <= "100110";
				when "0001110001011111" => data <= "100110";
				when "0001110001100000" => data <= "111111";
				when "0001110001101000" => data <= "111111";
				when "0001110001101001" => data <= "100110";
				when "0001110001101010" => data <= "100110";
				when "0001110001101011" => data <= "100110";
				when "0001110001101100" => data <= "100110";
				when "0001110001101101" => data <= "100110";
				when "0001110001101110" => data <= "100110";
				when "0001110001101111" => data <= "010110";
				when "0001110001110000" => data <= "100110";
				when "0001110001110001" => data <= "100110";
				when "0001110001110010" => data <= "010110";
				when "0001110001110011" => data <= "010110";
				when "0001110001110100" => data <= "111111";
				when "0001110100101000" => data <= "111111";
				when "0001110100101001" => data <= "010110";
				when "0001110100101010" => data <= "100110";
				when "0001110100101011" => data <= "100110";
				when "0001110100101100" => data <= "111111";
				when "0001110100111011" => data <= "111111";
				when "0001110100111100" => data <= "100110";
				when "0001110100111101" => data <= "100111";
				when "0001110100111110" => data <= "100111";
				when "0001110100111111" => data <= "100111";
				when "0001110101000000" => data <= "111111";
				when "0001110101000001" => data <= "111111";
				when "0001110101000010" => data <= "111111";
				when "0001110101000011" => data <= "100111";
				when "0001110101000100" => data <= "100111";
				when "0001110101000101" => data <= "100111";
				when "0001110101000110" => data <= "100110";
				when "0001110101000111" => data <= "111111";
				when "0001110101001111" => data <= "111111";
				when "0001110101010000" => data <= "100110";
				when "0001110101010001" => data <= "100111";
				when "0001110101010010" => data <= "100111";
				when "0001110101010011" => data <= "100111";
				when "0001110101010100" => data <= "100111";
				when "0001110101010101" => data <= "100110";
				when "0001110101010110" => data <= "111111";
				when "0001110101011001" => data <= "111111";
				when "0001110101011010" => data <= "100110";
				when "0001110101011011" => data <= "100110";
				when "0001110101011100" => data <= "100111";
				when "0001110101011101" => data <= "100111";
				when "0001110101011110" => data <= "100111";
				when "0001110101011111" => data <= "100110";
				when "0001110101100000" => data <= "111111";
				when "0001110101101000" => data <= "111111";
				when "0001110101101001" => data <= "100110";
				when "0001110101101010" => data <= "100111";
				when "0001110101101011" => data <= "100110";
				when "0001110101101100" => data <= "100110";
				when "0001110101101101" => data <= "111111";
				when "0001110101101110" => data <= "111111";
				when "0001110101101111" => data <= "111111";
				when "0001110101110000" => data <= "111111";
				when "0001110101110001" => data <= "111111";
				when "0001110101110010" => data <= "111111";
				when "0001110101110011" => data <= "111111";
				when "0001111000101000" => data <= "111111";
				when "0001111000101001" => data <= "100110";
				when "0001111000101010" => data <= "100110";
				when "0001111000101011" => data <= "100110";
				when "0001111000101100" => data <= "111111";
				when "0001111000111011" => data <= "111111";
				when "0001111000111100" => data <= "100110";
				when "0001111000111101" => data <= "100111";
				when "0001111000111110" => data <= "100110";
				when "0001111000111111" => data <= "100110";
				when "0001111001000000" => data <= "111111";
				when "0001111001000010" => data <= "111111";
				when "0001111001000011" => data <= "100111";
				when "0001111001000100" => data <= "100111";
				when "0001111001000101" => data <= "100111";
				when "0001111001000110" => data <= "100110";
				when "0001111001000111" => data <= "111111";
				when "0001111001001111" => data <= "111111";
				when "0001111001010000" => data <= "100110";
				when "0001111001010001" => data <= "100111";
				when "0001111001010010" => data <= "100111";
				when "0001111001010011" => data <= "100111";
				when "0001111001010100" => data <= "100111";
				when "0001111001010101" => data <= "100111";
				when "0001111001010110" => data <= "100110";
				when "0001111001010111" => data <= "111111";
				when "0001111001011000" => data <= "111111";
				when "0001111001011001" => data <= "100110";
				when "0001111001011010" => data <= "100111";
				when "0001111001011011" => data <= "100111";
				when "0001111001011100" => data <= "100111";
				when "0001111001011101" => data <= "100111";
				when "0001111001011110" => data <= "100111";
				when "0001111001011111" => data <= "100110";
				when "0001111001100000" => data <= "111111";
				when "0001111001101000" => data <= "111111";
				when "0001111001101001" => data <= "100110";
				when "0001111001101010" => data <= "100111";
				when "0001111001101011" => data <= "100110";
				when "0001111001101100" => data <= "100110";
				when "0001111001101101" => data <= "111111";
				when "0001111100101000" => data <= "111111";
				when "0001111100101001" => data <= "100110";
				when "0001111100101010" => data <= "100110";
				when "0001111100101011" => data <= "100110";
				when "0001111100101100" => data <= "111111";
				when "0001111100111011" => data <= "111111";
				when "0001111100111100" => data <= "100110";
				when "0001111100111101" => data <= "100111";
				when "0001111100111110" => data <= "100110";
				when "0001111100111111" => data <= "100110";
				when "0001111101000000" => data <= "111111";
				when "0001111101000001" => data <= "111111";
				when "0001111101000010" => data <= "111111";
				when "0001111101000011" => data <= "100111";
				when "0001111101000100" => data <= "100111";
				when "0001111101000101" => data <= "100111";
				when "0001111101000110" => data <= "100110";
				when "0001111101000111" => data <= "111111";
				when "0001111101001111" => data <= "111111";
				when "0001111101010000" => data <= "100110";
				when "0001111101010001" => data <= "100111";
				when "0001111101010010" => data <= "100111";
				when "0001111101010011" => data <= "100111";
				when "0001111101010100" => data <= "100111";
				when "0001111101010101" => data <= "100111";
				when "0001111101010110" => data <= "100111";
				when "0001111101010111" => data <= "100110";
				when "0001111101011000" => data <= "100110";
				when "0001111101011001" => data <= "100110";
				when "0001111101011010" => data <= "100111";
				when "0001111101011011" => data <= "100111";
				when "0001111101011100" => data <= "100111";
				when "0001111101011101" => data <= "100111";
				when "0001111101011110" => data <= "100111";
				when "0001111101011111" => data <= "100110";
				when "0001111101100000" => data <= "111111";
				when "0001111101101000" => data <= "111111";
				when "0001111101101001" => data <= "100110";
				when "0001111101101010" => data <= "100111";
				when "0001111101101011" => data <= "100110";
				when "0001111101101100" => data <= "100110";
				when "0001111101101101" => data <= "111111";
				when "0010000000101000" => data <= "111111";
				when "0010000000101001" => data <= "100110";
				when "0010000000101010" => data <= "100110";
				when "0010000000101011" => data <= "100110";
				when "0010000000101100" => data <= "111111";
				when "0010000000111011" => data <= "111111";
				when "0010000000111100" => data <= "100110";
				when "0010000000111101" => data <= "100111";
				when "0010000000111110" => data <= "100111";
				when "0010000000111111" => data <= "100111";
				when "0010000001000000" => data <= "100111";
				when "0010000001000001" => data <= "100110";
				when "0010000001000010" => data <= "100110";
				when "0010000001000011" => data <= "100111";
				when "0010000001000100" => data <= "100111";
				when "0010000001000101" => data <= "100111";
				when "0010000001000110" => data <= "100110";
				when "0010000001000111" => data <= "111111";
				when "0010000001001111" => data <= "111111";
				when "0010000001010000" => data <= "100110";
				when "0010000001010001" => data <= "100111";
				when "0010000001010010" => data <= "100110";
				when "0010000001010011" => data <= "100110";
				when "0010000001010100" => data <= "111111";
				when "0010000001010101" => data <= "100110";
				when "0010000001010110" => data <= "100111";
				when "0010000001010111" => data <= "100111";
				when "0010000001011000" => data <= "100111";
				when "0010000001011001" => data <= "100111";
				when "0010000001011010" => data <= "100110";
				when "0010000001011011" => data <= "111111";
				when "0010000001011100" => data <= "100111";
				when "0010000001011101" => data <= "100111";
				when "0010000001011110" => data <= "100111";
				when "0010000001011111" => data <= "100110";
				when "0010000001100000" => data <= "111111";
				when "0010000001101000" => data <= "111111";
				when "0010000001101001" => data <= "100111";
				when "0010000001101010" => data <= "100111";
				when "0010000001101011" => data <= "100110";
				when "0010000001101100" => data <= "100110";
				when "0010000001101101" => data <= "111111";
				when "0010000001101110" => data <= "111111";
				when "0010000001101111" => data <= "111111";
				when "0010000001110000" => data <= "111111";
				when "0010000001110001" => data <= "111111";
				when "0010000001110010" => data <= "111111";
				when "0010000001110011" => data <= "111111";
				when "0010000100101000" => data <= "111111";
				when "0010000100101001" => data <= "100110";
				when "0010000100101010" => data <= "100110";
				when "0010000100101011" => data <= "100110";
				when "0010000100101100" => data <= "111111";
				when "0010000100111011" => data <= "111111";
				when "0010000100111100" => data <= "100110";
				when "0010000100111101" => data <= "100111";
				when "0010000100111110" => data <= "100111";
				when "0010000100111111" => data <= "100111";
				when "0010000101000000" => data <= "100111";
				when "0010000101000001" => data <= "100110";
				when "0010000101000010" => data <= "100110";
				when "0010000101000011" => data <= "100111";
				when "0010000101000100" => data <= "100111";
				when "0010000101000101" => data <= "100111";
				when "0010000101000110" => data <= "100110";
				when "0010000101000111" => data <= "111111";
				when "0010000101001111" => data <= "111111";
				when "0010000101010000" => data <= "100110";
				when "0010000101010001" => data <= "100111";
				when "0010000101010010" => data <= "100110";
				when "0010000101010011" => data <= "100110";
				when "0010000101010100" => data <= "111111";
				when "0010000101010101" => data <= "100110";
				when "0010000101010110" => data <= "100111";
				when "0010000101010111" => data <= "100111";
				when "0010000101011000" => data <= "100111";
				when "0010000101011001" => data <= "100111";
				when "0010000101011010" => data <= "100110";
				when "0010000101011011" => data <= "111111";
				when "0010000101011100" => data <= "100111";
				when "0010000101011101" => data <= "100111";
				when "0010000101011110" => data <= "100111";
				when "0010000101011111" => data <= "100110";
				when "0010000101100000" => data <= "111111";
				when "0010000101101000" => data <= "111111";
				when "0010000101101001" => data <= "100111";
				when "0010000101101010" => data <= "100111";
				when "0010000101101011" => data <= "100110";
				when "0010000101101100" => data <= "100110";
				when "0010000101101101" => data <= "111111";
				when "0010000101101110" => data <= "111111";
				when "0010000101101111" => data <= "111111";
				when "0010000101110000" => data <= "111111";
				when "0010000101110001" => data <= "111111";
				when "0010000101110010" => data <= "111111";
				when "0010000101110011" => data <= "111111";
				when "0010001000101000" => data <= "111111";
				when "0010001000101001" => data <= "100110";
				when "0010001000101010" => data <= "100110";
				when "0010001000101011" => data <= "100110";
				when "0010001000101100" => data <= "111111";
				when "0010001000111011" => data <= "111111";
				when "0010001000111100" => data <= "100111";
				when "0010001000111101" => data <= "100111";
				when "0010001000111110" => data <= "100111";
				when "0010001000111111" => data <= "100111";
				when "0010001001000000" => data <= "100111";
				when "0010001001000001" => data <= "100110";
				when "0010001001000010" => data <= "100110";
				when "0010001001000011" => data <= "100111";
				when "0010001001000100" => data <= "100111";
				when "0010001001000101" => data <= "100111";
				when "0010001001000110" => data <= "100110";
				when "0010001001000111" => data <= "111111";
				when "0010001001001111" => data <= "111111";
				when "0010001001010000" => data <= "100110";
				when "0010001001010001" => data <= "100111";
				when "0010001001010010" => data <= "100110";
				when "0010001001010011" => data <= "100110";
				when "0010001001010100" => data <= "111111";
				when "0010001001010101" => data <= "111111";
				when "0010001001010110" => data <= "100110";
				when "0010001001010111" => data <= "100110";
				when "0010001001011000" => data <= "100110";
				when "0010001001011001" => data <= "100110";
				when "0010001001011010" => data <= "111111";
				when "0010001001011011" => data <= "111111";
				when "0010001001011100" => data <= "100111";
				when "0010001001011101" => data <= "100111";
				when "0010001001011110" => data <= "100111";
				when "0010001001011111" => data <= "100110";
				when "0010001001100000" => data <= "111111";
				when "0010001001101000" => data <= "111111";
				when "0010001001101001" => data <= "100111";
				when "0010001001101010" => data <= "100111";
				when "0010001001101011" => data <= "100111";
				when "0010001001101100" => data <= "100111";
				when "0010001001101101" => data <= "100110";
				when "0010001001101110" => data <= "100110";
				when "0010001001101111" => data <= "100110";
				when "0010001001110000" => data <= "100110";
				when "0010001001110001" => data <= "100110";
				when "0010001001110010" => data <= "100110";
				when "0010001001110011" => data <= "010110";
				when "0010001001110100" => data <= "111111";
				when "0010001100101000" => data <= "111111";
				when "0010001100101001" => data <= "010110";
				when "0010001100101010" => data <= "010010";
				when "0010001100101011" => data <= "010010";
				when "0010001100101100" => data <= "111111";
				when "0010001100111011" => data <= "111111";
				when "0010001100111100" => data <= "010010";
				when "0010001100111101" => data <= "010011";
				when "0010001100111110" => data <= "010010";
				when "0010001100111111" => data <= "010010";
				when "0010001101000000" => data <= "111111";
				when "0010001101000001" => data <= "111111";
				when "0010001101000010" => data <= "111111";
				when "0010001101000011" => data <= "010010";
				when "0010001101000100" => data <= "010010";
				when "0010001101000101" => data <= "010011";
				when "0010001101000110" => data <= "010010";
				when "0010001101000111" => data <= "111111";
				when "0010001101001111" => data <= "111111";
				when "0010001101010000" => data <= "010010";
				when "0010001101010001" => data <= "010010";
				when "0010001101010010" => data <= "010010";
				when "0010001101010011" => data <= "010010";
				when "0010001101010100" => data <= "111111";
				when "0010001101010101" => data <= "000001";
				when "0010001101010110" => data <= "111111";
				when "0010001101010111" => data <= "010110";
				when "0010001101011000" => data <= "010110";
				when "0010001101011001" => data <= "111111";
				when "0010001101011011" => data <= "111111";
				when "0010001101011100" => data <= "010010";
				when "0010001101011101" => data <= "010010";
				when "0010001101011110" => data <= "010010";
				when "0010001101011111" => data <= "010010";
				when "0010001101100000" => data <= "111111";
				when "0010001101101000" => data <= "111111";
				when "0010001101101001" => data <= "010010";
				when "0010001101101010" => data <= "010011";
				when "0010001101101011" => data <= "010010";
				when "0010001101101100" => data <= "010010";
				when "0010001101101101" => data <= "010010";
				when "0010001101101110" => data <= "010010";
				when "0010001101101111" => data <= "010010";
				when "0010001101110000" => data <= "010010";
				when "0010001101110001" => data <= "010010";
				when "0010001101110010" => data <= "010110";
				when "0010001101110011" => data <= "010101";
				when "0010001101110100" => data <= "111111";
				when "0010010000101000" => data <= "111111";
				when "0010010000101001" => data <= "010010";
				when "0010010000101010" => data <= "010110";
				when "0010010000101011" => data <= "010110";
				when "0010010000101100" => data <= "111111";
				when "0010010000111011" => data <= "111111";
				when "0010010000111100" => data <= "010010";
				when "0010010000111101" => data <= "010011";
				when "0010010000111110" => data <= "010010";
				when "0010010000111111" => data <= "010010";
				when "0010010001000000" => data <= "111111";
				when "0010010001000010" => data <= "111111";
				when "0010010001000011" => data <= "010010";
				when "0010010001000100" => data <= "010010";
				when "0010010001000101" => data <= "010011";
				when "0010010001000110" => data <= "010010";
				when "0010010001000111" => data <= "111111";
				when "0010010001001111" => data <= "111111";
				when "0010010001010000" => data <= "010010";
				when "0010010001010001" => data <= "010011";
				when "0010010001010010" => data <= "010010";
				when "0010010001010011" => data <= "010010";
				when "0010010001010100" => data <= "111111";
				when "0010010001010111" => data <= "111111";
				when "0010010001011000" => data <= "111111";
				when "0010010001011011" => data <= "111111";
				when "0010010001011100" => data <= "010010";
				when "0010010001011101" => data <= "010010";
				when "0010010001011110" => data <= "010011";
				when "0010010001011111" => data <= "010010";
				when "0010010001100000" => data <= "111111";
				when "0010010001101000" => data <= "111111";
				when "0010010001101001" => data <= "010010";
				when "0010010001101010" => data <= "010011";
				when "0010010001101011" => data <= "010010";
				when "0010010001101100" => data <= "010010";
				when "0010010001101101" => data <= "111111";
				when "0010010001101110" => data <= "111111";
				when "0010010001101111" => data <= "111111";
				when "0010010001110000" => data <= "111111";
				when "0010010001110001" => data <= "111111";
				when "0010010001110010" => data <= "111111";
				when "0010010001110011" => data <= "111111";
				when "0010010100101000" => data <= "111111";
				when "0010010100101001" => data <= "010110";
				when "0010010100101010" => data <= "010110";
				when "0010010100101011" => data <= "010110";
				when "0010010100101100" => data <= "111111";
				when "0010010100101110" => data <= "111111";
				when "0010010100101111" => data <= "111111";
				when "0010010100110000" => data <= "111111";
				when "0010010100110001" => data <= "111111";
				when "0010010100110010" => data <= "111111";
				when "0010010100110011" => data <= "111111";
				when "0010010100111011" => data <= "111111";
				when "0010010100111100" => data <= "010010";
				when "0010010100111101" => data <= "010011";
				when "0010010100111110" => data <= "010010";
				when "0010010100111111" => data <= "010010";
				when "0010010101000000" => data <= "111111";
				when "0010010101000010" => data <= "111111";
				when "0010010101000011" => data <= "010010";
				when "0010010101000100" => data <= "010010";
				when "0010010101000101" => data <= "010011";
				when "0010010101000110" => data <= "010010";
				when "0010010101000111" => data <= "111111";
				when "0010010101001111" => data <= "111111";
				when "0010010101010000" => data <= "010010";
				when "0010010101010001" => data <= "010011";
				when "0010010101010010" => data <= "010010";
				when "0010010101010011" => data <= "010010";
				when "0010010101010100" => data <= "111111";
				when "0010010101011011" => data <= "111111";
				when "0010010101011100" => data <= "010010";
				when "0010010101011101" => data <= "010010";
				when "0010010101011110" => data <= "010011";
				when "0010010101011111" => data <= "010010";
				when "0010010101100000" => data <= "111111";
				when "0010010101101000" => data <= "111111";
				when "0010010101101001" => data <= "010010";
				when "0010010101101010" => data <= "010011";
				when "0010010101101011" => data <= "010010";
				when "0010010101101100" => data <= "010010";
				when "0010010101101101" => data <= "111111";
				when "0010010101101110" => data <= "000001";
				when "0010011000101000" => data <= "111111";
				when "0010011000101001" => data <= "010110";
				when "0010011000101010" => data <= "010110";
				when "0010011000101011" => data <= "010110";
				when "0010011000101100" => data <= "111111";
				when "0010011000101110" => data <= "111111";
				when "0010011000101111" => data <= "111111";
				when "0010011000110000" => data <= "111111";
				when "0010011000110001" => data <= "111111";
				when "0010011000110010" => data <= "111111";
				when "0010011000110011" => data <= "111111";
				when "0010011000111011" => data <= "111111";
				when "0010011000111100" => data <= "010010";
				when "0010011000111101" => data <= "010011";
				when "0010011000111110" => data <= "010010";
				when "0010011000111111" => data <= "010010";
				when "0010011001000000" => data <= "111111";
				when "0010011001000010" => data <= "111111";
				when "0010011001000011" => data <= "010010";
				when "0010011001000100" => data <= "010010";
				when "0010011001000101" => data <= "010011";
				when "0010011001000110" => data <= "010010";
				when "0010011001000111" => data <= "111111";
				when "0010011001001111" => data <= "111111";
				when "0010011001010000" => data <= "010010";
				when "0010011001010001" => data <= "010011";
				when "0010011001010010" => data <= "010010";
				when "0010011001010011" => data <= "010010";
				when "0010011001010100" => data <= "111111";
				when "0010011001011011" => data <= "111111";
				when "0010011001011100" => data <= "010010";
				when "0010011001011101" => data <= "010010";
				when "0010011001011110" => data <= "010011";
				when "0010011001011111" => data <= "010010";
				when "0010011001100000" => data <= "111111";
				when "0010011001101000" => data <= "111111";
				when "0010011001101001" => data <= "010010";
				when "0010011001101010" => data <= "010011";
				when "0010011001101011" => data <= "010010";
				when "0010011001101100" => data <= "010010";
				when "0010011001101101" => data <= "111111";
				when "0010011001101110" => data <= "000001";
				when "0010011100101000" => data <= "111111";
				when "0010011100101001" => data <= "010110";
				when "0010011100101010" => data <= "010010";
				when "0010011100101011" => data <= "010010";
				when "0010011100101100" => data <= "111111";
				when "0010011100101110" => data <= "111111";
				when "0010011100101111" => data <= "010001";
				when "0010011100110000" => data <= "010001";
				when "0010011100110001" => data <= "010001";
				when "0010011100110010" => data <= "010001";
				when "0010011100110011" => data <= "111111";
				when "0010011100111011" => data <= "111111";
				when "0010011100111100" => data <= "010010";
				when "0010011100111101" => data <= "010010";
				when "0010011100111110" => data <= "010010";
				when "0010011100111111" => data <= "010010";
				when "0010011101000000" => data <= "111111";
				when "0010011101000010" => data <= "111111";
				when "0010011101000011" => data <= "010010";
				when "0010011101000100" => data <= "010010";
				when "0010011101000101" => data <= "010011";
				when "0010011101000110" => data <= "010010";
				when "0010011101000111" => data <= "111111";
				when "0010011101001111" => data <= "111111";
				when "0010011101010000" => data <= "010010";
				when "0010011101010001" => data <= "010011";
				when "0010011101010010" => data <= "010010";
				when "0010011101010011" => data <= "010010";
				when "0010011101010100" => data <= "111111";
				when "0010011101011011" => data <= "111111";
				when "0010011101011100" => data <= "010010";
				when "0010011101011101" => data <= "010010";
				when "0010011101011110" => data <= "010011";
				when "0010011101011111" => data <= "010110";
				when "0010011101100000" => data <= "111111";
				when "0010011101101000" => data <= "111111";
				when "0010011101101001" => data <= "010010";
				when "0010011101101010" => data <= "010011";
				when "0010011101101011" => data <= "010010";
				when "0010011101101100" => data <= "010010";
				when "0010011101101101" => data <= "111111";
				when "0010100000101000" => data <= "111111";
				when "0010100000101001" => data <= "010110";
				when "0010100000101010" => data <= "010110";
				when "0010100000101011" => data <= "010110";
				when "0010100000101100" => data <= "111111";
				when "0010100000101110" => data <= "111111";
				when "0010100000101111" => data <= "111111";
				when "0010100000110000" => data <= "111111";
				when "0010100000110001" => data <= "010001";
				when "0010100000110010" => data <= "010001";
				when "0010100000110011" => data <= "111111";
				when "0010100000111011" => data <= "111111";
				when "0010100000111100" => data <= "010010";
				when "0010100000111101" => data <= "010010";
				when "0010100000111110" => data <= "010010";
				when "0010100000111111" => data <= "010010";
				when "0010100001000000" => data <= "111111";
				when "0010100001000010" => data <= "111111";
				when "0010100001000011" => data <= "010010";
				when "0010100001000100" => data <= "010010";
				when "0010100001000101" => data <= "010010";
				when "0010100001000110" => data <= "010010";
				when "0010100001000111" => data <= "111111";
				when "0010100001001111" => data <= "111111";
				when "0010100001010000" => data <= "010010";
				when "0010100001010001" => data <= "010010";
				when "0010100001010010" => data <= "010010";
				when "0010100001010011" => data <= "010010";
				when "0010100001010100" => data <= "111111";
				when "0010100001011011" => data <= "111111";
				when "0010100001011100" => data <= "010010";
				when "0010100001011101" => data <= "010010";
				when "0010100001011110" => data <= "010010";
				when "0010100001011111" => data <= "010010";
				when "0010100001100000" => data <= "111111";
				when "0010100001101000" => data <= "111111";
				when "0010100001101001" => data <= "010010";
				when "0010100001101010" => data <= "010010";
				when "0010100001101011" => data <= "010010";
				when "0010100001101100" => data <= "010010";
				when "0010100001101101" => data <= "111111";
				when "0010100100101000" => data <= "111111";
				when "0010100100101001" => data <= "010001";
				when "0010100100101010" => data <= "000001";
				when "0010100100101011" => data <= "000001";
				when "0010100100101100" => data <= "111111";
				when "0010100100101101" => data <= "000001";
				when "0010100100101110" => data <= "000001";
				when "0010100100101111" => data <= "111111";
				when "0010100100110000" => data <= "111111";
				when "0010100100110001" => data <= "000001";
				when "0010100100110010" => data <= "010001";
				when "0010100100110011" => data <= "111111";
				when "0010100100111011" => data <= "111111";
				when "0010100100111100" => data <= "010010";
				when "0010100100111101" => data <= "010010";
				when "0010100100111110" => data <= "010010";
				when "0010100100111111" => data <= "010010";
				when "0010100101000000" => data <= "111111";
				when "0010100101000010" => data <= "111111";
				when "0010100101000011" => data <= "010010";
				when "0010100101000100" => data <= "010010";
				when "0010100101000101" => data <= "010010";
				when "0010100101000110" => data <= "010010";
				when "0010100101000111" => data <= "111111";
				when "0010100101001111" => data <= "111111";
				when "0010100101010000" => data <= "010010";
				when "0010100101010001" => data <= "000010";
				when "0010100101010010" => data <= "010010";
				when "0010100101010011" => data <= "010010";
				when "0010100101010100" => data <= "111111";
				when "0010100101011011" => data <= "111111";
				when "0010100101011100" => data <= "000010";
				when "0010100101011101" => data <= "000010";
				when "0010100101011110" => data <= "010010";
				when "0010100101011111" => data <= "000010";
				when "0010100101100000" => data <= "111111";
				when "0010100101101000" => data <= "111111";
				when "0010100101101001" => data <= "010010";
				when "0010100101101010" => data <= "010010";
				when "0010100101101011" => data <= "010010";
				when "0010100101101100" => data <= "010010";
				when "0010100101101101" => data <= "111111";
				when "0010100101101110" => data <= "111111";
				when "0010100101101111" => data <= "111111";
				when "0010100101110000" => data <= "111111";
				when "0010100101110001" => data <= "111111";
				when "0010100101110010" => data <= "111111";
				when "0010100101110011" => data <= "111111";
				when "0010101000101000" => data <= "111111";
				when "0010101000101001" => data <= "010001";
				when "0010101000101010" => data <= "000010";
				when "0010101000101011" => data <= "000010";
				when "0010101000101100" => data <= "111111";
				when "0010101000101101" => data <= "111111";
				when "0010101000101110" => data <= "111111";
				when "0010101000101111" => data <= "111111";
				when "0010101000110000" => data <= "111111";
				when "0010101000110001" => data <= "010010";
				when "0010101000110010" => data <= "010001";
				when "0010101000110011" => data <= "111111";
				when "0010101000111011" => data <= "111111";
				when "0010101000111100" => data <= "010010";
				when "0010101000111101" => data <= "010010";
				when "0010101000111110" => data <= "010010";
				when "0010101000111111" => data <= "010010";
				when "0010101001000000" => data <= "111111";
				when "0010101001000010" => data <= "111111";
				when "0010101001000011" => data <= "010010";
				when "0010101001000100" => data <= "010010";
				when "0010101001000101" => data <= "010010";
				when "0010101001000110" => data <= "010010";
				when "0010101001000111" => data <= "111111";
				when "0010101001001111" => data <= "111111";
				when "0010101001010000" => data <= "000010";
				when "0010101001010001" => data <= "010010";
				when "0010101001010010" => data <= "000010";
				when "0010101001010011" => data <= "000010";
				when "0010101001010100" => data <= "111111";
				when "0010101001011011" => data <= "111111";
				when "0010101001011100" => data <= "000010";
				when "0010101001011101" => data <= "000010";
				when "0010101001011110" => data <= "000010";
				when "0010101001011111" => data <= "010010";
				when "0010101001100000" => data <= "111111";
				when "0010101001101000" => data <= "111111";
				when "0010101001101001" => data <= "010010";
				when "0010101001101010" => data <= "010010";
				when "0010101001101011" => data <= "000010";
				when "0010101001101100" => data <= "000010";
				when "0010101001101101" => data <= "000010";
				when "0010101001101110" => data <= "010010";
				when "0010101001101111" => data <= "010010";
				when "0010101001110000" => data <= "010010";
				when "0010101001110001" => data <= "010010";
				when "0010101001110010" => data <= "010010";
				when "0010101001110011" => data <= "000001";
				when "0010101001110100" => data <= "111111";
				when "0010101100101000" => data <= "111111";
				when "0010101100101001" => data <= "010001";
				when "0010101100101010" => data <= "000010";
				when "0010101100101011" => data <= "000010";
				when "0010101100101100" => data <= "111111";
				when "0010101100101101" => data <= "111111";
				when "0010101100101110" => data <= "111111";
				when "0010101100101111" => data <= "111111";
				when "0010101100110000" => data <= "111111";
				when "0010101100110001" => data <= "010010";
				when "0010101100110010" => data <= "010001";
				when "0010101100110011" => data <= "111111";
				when "0010101100111011" => data <= "111111";
				when "0010101100111100" => data <= "010010";
				when "0010101100111101" => data <= "010010";
				when "0010101100111110" => data <= "010010";
				when "0010101100111111" => data <= "010010";
				when "0010101101000000" => data <= "111111";
				when "0010101101000010" => data <= "111111";
				when "0010101101000011" => data <= "010010";
				when "0010101101000100" => data <= "010010";
				when "0010101101000101" => data <= "010010";
				when "0010101101000110" => data <= "010010";
				when "0010101101000111" => data <= "111111";
				when "0010101101001111" => data <= "111111";
				when "0010101101010000" => data <= "000010";
				when "0010101101010001" => data <= "010010";
				when "0010101101010010" => data <= "000010";
				when "0010101101010011" => data <= "000010";
				when "0010101101010100" => data <= "111111";
				when "0010101101011011" => data <= "111111";
				when "0010101101011100" => data <= "000010";
				when "0010101101011101" => data <= "000010";
				when "0010101101011110" => data <= "000010";
				when "0010101101011111" => data <= "010010";
				when "0010101101100000" => data <= "111111";
				when "0010101101101000" => data <= "111111";
				when "0010101101101001" => data <= "010010";
				when "0010101101101010" => data <= "010010";
				when "0010101101101011" => data <= "000010";
				when "0010101101101100" => data <= "000010";
				when "0010101101101101" => data <= "000010";
				when "0010101101101110" => data <= "010010";
				when "0010101101101111" => data <= "010010";
				when "0010101101110000" => data <= "010010";
				when "0010101101110001" => data <= "010010";
				when "0010101101110010" => data <= "010010";
				when "0010101101110011" => data <= "000001";
				when "0010101101110100" => data <= "111111";
				when "0010110000101000" => data <= "111111";
				when "0010110000101001" => data <= "000001";
				when "0010110000101010" => data <= "010001";
				when "0010110000101011" => data <= "010001";
				when "0010110000101100" => data <= "010001";
				when "0010110000101101" => data <= "010001";
				when "0010110000101110" => data <= "010001";
				when "0010110000101111" => data <= "010001";
				when "0010110000110000" => data <= "010001";
				when "0010110000110001" => data <= "000001";
				when "0010110000110010" => data <= "000001";
				when "0010110000110011" => data <= "111111";
				when "0010110000111011" => data <= "111111";
				when "0010110000111100" => data <= "010010";
				when "0010110000111101" => data <= "010010";
				when "0010110000111110" => data <= "010001";
				when "0010110000111111" => data <= "010001";
				when "0010110001000000" => data <= "111111";
				when "0010110001000010" => data <= "111111";
				when "0010110001000011" => data <= "010001";
				when "0010110001000100" => data <= "010001";
				when "0010110001000101" => data <= "010010";
				when "0010110001000110" => data <= "010001";
				when "0010110001000111" => data <= "111111";
				when "0010110001001111" => data <= "111111";
				when "0010110001010000" => data <= "000001";
				when "0010110001010001" => data <= "000010";
				when "0010110001010010" => data <= "000001";
				when "0010110001010011" => data <= "000001";
				when "0010110001010100" => data <= "111111";
				when "0010110001011011" => data <= "111111";
				when "0010110001011100" => data <= "000001";
				when "0010110001011101" => data <= "000001";
				when "0010110001011110" => data <= "010010";
				when "0010110001011111" => data <= "000001";
				when "0010110001100000" => data <= "111111";
				when "0010110001101000" => data <= "111111";
				when "0010110001101001" => data <= "010010";
				when "0010110001101010" => data <= "000010";
				when "0010110001101011" => data <= "010010";
				when "0010110001101100" => data <= "010010";
				when "0010110001101101" => data <= "000010";
				when "0010110001101110" => data <= "010010";
				when "0010110001101111" => data <= "010010";
				when "0010110001110000" => data <= "010010";
				when "0010110001110001" => data <= "010010";
				when "0010110001110010" => data <= "010010";
				when "0010110001110011" => data <= "000001";
				when "0010110001110100" => data <= "111111";
				when "0010110100101001" => data <= "111111";
				when "0010110100101010" => data <= "111111";
				when "0010110100101011" => data <= "111111";
				when "0010110100101100" => data <= "111111";
				when "0010110100101101" => data <= "111111";
				when "0010110100101110" => data <= "111111";
				when "0010110100101111" => data <= "111111";
				when "0010110100110000" => data <= "111111";
				when "0010110100110001" => data <= "111111";
				when "0010110100110010" => data <= "111111";
				when "0010110100111100" => data <= "111111";
				when "0010110100111101" => data <= "111111";
				when "0010110100111110" => data <= "111111";
				when "0010110100111111" => data <= "111111";
				when "0010110101000011" => data <= "111111";
				when "0010110101000100" => data <= "111111";
				when "0010110101000101" => data <= "111111";
				when "0010110101000110" => data <= "111111";
				when "0010110101010000" => data <= "111111";
				when "0010110101010001" => data <= "111111";
				when "0010110101010010" => data <= "111111";
				when "0010110101010011" => data <= "111111";
				when "0010110101011100" => data <= "111111";
				when "0010110101011101" => data <= "111111";
				when "0010110101011110" => data <= "111111";
				when "0010110101011111" => data <= "111111";
				when "0010110101101010" => data <= "111111";
				when "0010110101101011" => data <= "111111";
				when "0010110101101100" => data <= "111111";
				when "0010110101101101" => data <= "111111";
				when "0010110101101110" => data <= "111111";
				when "0010110101101111" => data <= "111111";
				when "0010110101110000" => data <= "111111";
				when "0010110101110001" => data <= "111111";
				when "0010110101110010" => data <= "111111";
				when "0010110101110011" => data <= "111111";
				when "0011010000101000" => data <= "111111";
				when "0011010000101001" => data <= "111111";
				when "0011010000101010" => data <= "111111";
				when "0011010000101011" => data <= "111111";
				when "0011010000101100" => data <= "111111";
				when "0011010000101101" => data <= "111111";
				when "0011010000101110" => data <= "111111";
				when "0011010000101111" => data <= "111111";
				when "0011010000110000" => data <= "111111";
				when "0011010000110001" => data <= "111111";
				when "0011010000110010" => data <= "111111";
				when "0011010000110011" => data <= "111111";
				when "0011010000111011" => data <= "111111";
				when "0011010000111100" => data <= "111111";
				when "0011010000111101" => data <= "111111";
				when "0011010000111110" => data <= "111111";
				when "0011010000111111" => data <= "111111";
				when "0011010001000000" => data <= "111111";
				when "0011010001001010" => data <= "111111";
				when "0011010001001011" => data <= "111111";
				when "0011010001001100" => data <= "111111";
				when "0011010001001101" => data <= "111111";
				when "0011010001001110" => data <= "111111";
				when "0011010001001111" => data <= "111111";
				when "0011010001010111" => data <= "111111";
				when "0011010001011000" => data <= "111111";
				when "0011010001011001" => data <= "111111";
				when "0011010001011010" => data <= "111111";
				when "0011010001011011" => data <= "111111";
				when "0011010001011100" => data <= "111111";
				when "0011010001011101" => data <= "111111";
				when "0011010001011110" => data <= "111111";
				when "0011010001011111" => data <= "111111";
				when "0011010001100000" => data <= "111111";
				when "0011010001100001" => data <= "111111";
				when "0011010001100010" => data <= "111111";
				when "0011010001101010" => data <= "111111";
				when "0011010001101011" => data <= "111111";
				when "0011010001101100" => data <= "111111";
				when "0011010001101101" => data <= "111111";
				when "0011010001101110" => data <= "111111";
				when "0011010001101111" => data <= "111111";
				when "0011010001110000" => data <= "111111";
				when "0011010001110001" => data <= "111111";
				when "0011010001110010" => data <= "111111";
				when "0011010001110011" => data <= "111111";
				when "0011010001110100" => data <= "111111";
				when "0011010100101000" => data <= "111111";
				when "0011010100101001" => data <= "111111";
				when "0011010100101010" => data <= "111111";
				when "0011010100101011" => data <= "111111";
				when "0011010100101100" => data <= "111111";
				when "0011010100101101" => data <= "111111";
				when "0011010100101110" => data <= "111111";
				when "0011010100101111" => data <= "111111";
				when "0011010100110000" => data <= "111111";
				when "0011010100110001" => data <= "111111";
				when "0011010100110010" => data <= "111111";
				when "0011010100110011" => data <= "111111";
				when "0011010100111011" => data <= "111111";
				when "0011010100111100" => data <= "111111";
				when "0011010100111101" => data <= "111111";
				when "0011010100111110" => data <= "111111";
				when "0011010100111111" => data <= "111111";
				when "0011010101000000" => data <= "111111";
				when "0011010101001010" => data <= "111111";
				when "0011010101001011" => data <= "111111";
				when "0011010101001100" => data <= "111111";
				when "0011010101001101" => data <= "111111";
				when "0011010101001110" => data <= "111111";
				when "0011010101001111" => data <= "111111";
				when "0011010101010111" => data <= "111111";
				when "0011010101011000" => data <= "111111";
				when "0011010101011001" => data <= "111111";
				when "0011010101011010" => data <= "111111";
				when "0011010101011011" => data <= "111111";
				when "0011010101011100" => data <= "111111";
				when "0011010101011101" => data <= "111111";
				when "0011010101011110" => data <= "111111";
				when "0011010101011111" => data <= "111111";
				when "0011010101100000" => data <= "111111";
				when "0011010101100001" => data <= "111111";
				when "0011010101100010" => data <= "111111";
				when "0011010101101010" => data <= "111111";
				when "0011010101101011" => data <= "111111";
				when "0011010101101100" => data <= "111111";
				when "0011010101101101" => data <= "111111";
				when "0011010101101110" => data <= "111111";
				when "0011010101101111" => data <= "111111";
				when "0011010101110000" => data <= "111111";
				when "0011010101110001" => data <= "111111";
				when "0011010101110010" => data <= "111111";
				when "0011010101110011" => data <= "111111";
				when "0011010101110100" => data <= "111111";
				when "0011011000100111" => data <= "111111";
				when "0011011000101000" => data <= "100110";
				when "0011011000101001" => data <= "100110";
				when "0011011000101010" => data <= "100110";
				when "0011011000101011" => data <= "100110";
				when "0011011000101100" => data <= "100110";
				when "0011011000101101" => data <= "100110";
				when "0011011000101110" => data <= "100110";
				when "0011011000101111" => data <= "100110";
				when "0011011000110000" => data <= "100110";
				when "0011011000110001" => data <= "100110";
				when "0011011000110010" => data <= "100110";
				when "0011011000110011" => data <= "010110";
				when "0011011000110100" => data <= "111111";
				when "0011011000110101" => data <= "111111";
				when "0011011000111011" => data <= "111111";
				when "0011011000111100" => data <= "100110";
				when "0011011000111101" => data <= "100110";
				when "0011011000111110" => data <= "100110";
				when "0011011000111111" => data <= "100110";
				when "0011011001000000" => data <= "111111";
				when "0011011001001010" => data <= "111111";
				when "0011011001001011" => data <= "010110";
				when "0011011001001100" => data <= "100110";
				when "0011011001001101" => data <= "010110";
				when "0011011001001110" => data <= "010110";
				when "0011011001001111" => data <= "111111";
				when "0011011001010110" => data <= "111111";
				when "0011011001010111" => data <= "100110";
				when "0011011001011000" => data <= "100110";
				when "0011011001011001" => data <= "100110";
				when "0011011001011010" => data <= "100110";
				when "0011011001011011" => data <= "100110";
				when "0011011001011100" => data <= "100110";
				when "0011011001011101" => data <= "100110";
				when "0011011001011110" => data <= "010110";
				when "0011011001011111" => data <= "100110";
				when "0011011001100000" => data <= "100110";
				when "0011011001100001" => data <= "010110";
				when "0011011001100010" => data <= "010110";
				when "0011011001100011" => data <= "111111";
				when "0011011001101001" => data <= "111111";
				when "0011011001101010" => data <= "010110";
				when "0011011001101011" => data <= "100110";
				when "0011011001101100" => data <= "100110";
				when "0011011001101101" => data <= "100110";
				when "0011011001101110" => data <= "100110";
				when "0011011001101111" => data <= "010110";
				when "0011011001110000" => data <= "100110";
				when "0011011001110001" => data <= "100110";
				when "0011011001110010" => data <= "100110";
				when "0011011001110011" => data <= "100110";
				when "0011011001110100" => data <= "100110";
				when "0011011001110101" => data <= "111111";
				when "0011011001110110" => data <= "111111";
				when "0011011100100111" => data <= "111111";
				when "0011011100101000" => data <= "100110";
				when "0011011100101001" => data <= "100110";
				when "0011011100101010" => data <= "100110";
				when "0011011100101011" => data <= "100110";
				when "0011011100101100" => data <= "100110";
				when "0011011100101101" => data <= "100110";
				when "0011011100101110" => data <= "100110";
				when "0011011100101111" => data <= "100110";
				when "0011011100110000" => data <= "100110";
				when "0011011100110001" => data <= "100110";
				when "0011011100110010" => data <= "100110";
				when "0011011100110011" => data <= "100110";
				when "0011011100110100" => data <= "111111";
				when "0011011100110101" => data <= "111111";
				when "0011011100111011" => data <= "111111";
				when "0011011100111100" => data <= "100110";
				when "0011011100111101" => data <= "100111";
				when "0011011100111110" => data <= "100110";
				when "0011011100111111" => data <= "100110";
				when "0011011101000000" => data <= "111011";
				when "0011011101000001" => data <= "111111";
				when "0011011101001000" => data <= "111111";
				when "0011011101001001" => data <= "111111";
				when "0011011101001010" => data <= "111111";
				when "0011011101001011" => data <= "100110";
				when "0011011101001100" => data <= "100110";
				when "0011011101001101" => data <= "100110";
				when "0011011101001110" => data <= "100110";
				when "0011011101001111" => data <= "111111";
				when "0011011101010110" => data <= "111111";
				when "0011011101010111" => data <= "010110";
				when "0011011101011000" => data <= "010110";
				when "0011011101011001" => data <= "100111";
				when "0011011101011010" => data <= "100110";
				when "0011011101011011" => data <= "100110";
				when "0011011101011100" => data <= "100110";
				when "0011011101011101" => data <= "100110";
				when "0011011101011110" => data <= "010110";
				when "0011011101011111" => data <= "100110";
				when "0011011101100000" => data <= "010110";
				when "0011011101100001" => data <= "010110";
				when "0011011101100010" => data <= "010110";
				when "0011011101100011" => data <= "111111";
				when "0011011101101001" => data <= "111111";
				when "0011011101101010" => data <= "100110";
				when "0011011101101011" => data <= "100110";
				when "0011011101101100" => data <= "100110";
				when "0011011101101101" => data <= "100110";
				when "0011011101101110" => data <= "100110";
				when "0011011101101111" => data <= "100110";
				when "0011011101110000" => data <= "100110";
				when "0011011101110001" => data <= "100110";
				when "0011011101110010" => data <= "100110";
				when "0011011101110011" => data <= "100111";
				when "0011011101110100" => data <= "100110";
				when "0011011101110101" => data <= "111111";
				when "0011011101110110" => data <= "111111";
				when "0011100000100111" => data <= "111111";
				when "0011100000101000" => data <= "100110";
				when "0011100000101001" => data <= "100110";
				when "0011100000101010" => data <= "111111";
				when "0011100000101011" => data <= "111111";
				when "0011100000101100" => data <= "111111";
				when "0011100000101101" => data <= "111111";
				when "0011100000101110" => data <= "111111";
				when "0011100000101111" => data <= "111111";
				when "0011100000110000" => data <= "111111";
				when "0011100000110001" => data <= "111111";
				when "0011100000110010" => data <= "100111";
				when "0011100000110011" => data <= "100111";
				when "0011100000110100" => data <= "111111";
				when "0011100000110101" => data <= "111111";
				when "0011100000111011" => data <= "111111";
				when "0011100000111100" => data <= "100110";
				when "0011100000111101" => data <= "100111";
				when "0011100000111110" => data <= "100110";
				when "0011100000111111" => data <= "100110";
				when "0011100001000000" => data <= "100110";
				when "0011100001000001" => data <= "111111";
				when "0011100001001000" => data <= "111111";
				when "0011100001001001" => data <= "111111";
				when "0011100001001010" => data <= "100110";
				when "0011100001001011" => data <= "100111";
				when "0011100001001100" => data <= "100111";
				when "0011100001001101" => data <= "100110";
				when "0011100001001110" => data <= "100110";
				when "0011100001001111" => data <= "111111";
				when "0011100001010110" => data <= "111111";
				when "0011100001010111" => data <= "100110";
				when "0011100001011000" => data <= "100110";
				when "0011100001011001" => data <= "100111";
				when "0011100001011010" => data <= "100110";
				when "0011100001011011" => data <= "111111";
				when "0011100001011100" => data <= "111111";
				when "0011100001011101" => data <= "111111";
				when "0011100001011110" => data <= "111111";
				when "0011100001011111" => data <= "111111";
				when "0011100001100000" => data <= "111111";
				when "0011100001100001" => data <= "111111";
				when "0011100001100010" => data <= "111111";
				when "0011100001101001" => data <= "111111";
				when "0011100001101010" => data <= "100110";
				when "0011100001101011" => data <= "100111";
				when "0011100001101100" => data <= "100111";
				when "0011100001101101" => data <= "100111";
				when "0011100001101110" => data <= "111111";
				when "0011100001101111" => data <= "111111";
				when "0011100001110000" => data <= "111111";
				when "0011100001110001" => data <= "111111";
				when "0011100001110010" => data <= "100110";
				when "0011100001110011" => data <= "100111";
				when "0011100001110100" => data <= "100110";
				when "0011100001110101" => data <= "111111";
				when "0011100001110110" => data <= "111111";
				when "0011100100100111" => data <= "111111";
				when "0011100100101000" => data <= "100110";
				when "0011100100101001" => data <= "100110";
				when "0011100100101010" => data <= "111111";
				when "0011100100101011" => data <= "111111";
				when "0011100100110001" => data <= "111111";
				when "0011100100110010" => data <= "100110";
				when "0011100100110011" => data <= "100110";
				when "0011100100110100" => data <= "111111";
				when "0011100100110101" => data <= "111111";
				when "0011100100111011" => data <= "111111";
				when "0011100100111100" => data <= "111111";
				when "0011100100111101" => data <= "100110";
				when "0011100100111110" => data <= "100110";
				when "0011100100111111" => data <= "100110";
				when "0011100101000000" => data <= "100110";
				when "0011100101000001" => data <= "111111";
				when "0011100101000111" => data <= "111111";
				when "0011100101001000" => data <= "111111";
				when "0011100101001001" => data <= "111111";
				when "0011100101001010" => data <= "010110";
				when "0011100101001011" => data <= "100110";
				when "0011100101001100" => data <= "100110";
				when "0011100101001101" => data <= "111111";
				when "0011100101001110" => data <= "111111";
				when "0011100101001111" => data <= "111111";
				when "0011100101010110" => data <= "111111";
				when "0011100101010111" => data <= "100110";
				when "0011100101011000" => data <= "100110";
				when "0011100101011001" => data <= "100111";
				when "0011100101011010" => data <= "100110";
				when "0011100101011011" => data <= "111111";
				when "0011100101101001" => data <= "111111";
				when "0011100101101010" => data <= "100110";
				when "0011100101101011" => data <= "100111";
				when "0011100101101100" => data <= "100111";
				when "0011100101101101" => data <= "100110";
				when "0011100101101110" => data <= "111111";
				when "0011100101110010" => data <= "111111";
				when "0011100101110011" => data <= "100111";
				when "0011100101110100" => data <= "100110";
				when "0011100101110101" => data <= "111111";
				when "0011100101110110" => data <= "111111";
				when "0011101000100111" => data <= "111111";
				when "0011101000101000" => data <= "100110";
				when "0011101000101001" => data <= "100110";
				when "0011101000101010" => data <= "111111";
				when "0011101000101011" => data <= "111111";
				when "0011101000110001" => data <= "111111";
				when "0011101000110010" => data <= "100110";
				when "0011101000110011" => data <= "100110";
				when "0011101000110100" => data <= "111111";
				when "0011101000110101" => data <= "111111";
				when "0011101000111011" => data <= "111111";
				when "0011101000111100" => data <= "111111";
				when "0011101000111101" => data <= "100110";
				when "0011101000111110" => data <= "100110";
				when "0011101000111111" => data <= "100110";
				when "0011101001000000" => data <= "100110";
				when "0011101001000001" => data <= "111111";
				when "0011101001000111" => data <= "111111";
				when "0011101001001000" => data <= "111111";
				when "0011101001001001" => data <= "111111";
				when "0011101001001010" => data <= "010110";
				when "0011101001001011" => data <= "100110";
				when "0011101001001100" => data <= "100110";
				when "0011101001001101" => data <= "111111";
				when "0011101001001110" => data <= "111111";
				when "0011101001001111" => data <= "111111";
				when "0011101001010110" => data <= "111111";
				when "0011101001010111" => data <= "100110";
				when "0011101001011000" => data <= "100110";
				when "0011101001011001" => data <= "100111";
				when "0011101001011010" => data <= "100110";
				when "0011101001011011" => data <= "111111";
				when "0011101001101001" => data <= "111111";
				when "0011101001101010" => data <= "100110";
				when "0011101001101011" => data <= "100111";
				when "0011101001101100" => data <= "100111";
				when "0011101001101101" => data <= "100110";
				when "0011101001101110" => data <= "111111";
				when "0011101001110010" => data <= "111111";
				when "0011101001110011" => data <= "100111";
				when "0011101001110100" => data <= "100110";
				when "0011101001110101" => data <= "111111";
				when "0011101001110110" => data <= "111111";
				when "0011101100100111" => data <= "111111";
				when "0011101100101000" => data <= "100111";
				when "0011101100101001" => data <= "100111";
				when "0011101100101010" => data <= "111111";
				when "0011101100101011" => data <= "111111";
				when "0011101100110001" => data <= "111111";
				when "0011101100110010" => data <= "100111";
				when "0011101100110011" => data <= "100110";
				when "0011101100110100" => data <= "111111";
				when "0011101100110101" => data <= "111111";
				when "0011101100111100" => data <= "111111";
				when "0011101100111101" => data <= "010110";
				when "0011101100111110" => data <= "100111";
				when "0011101100111111" => data <= "100111";
				when "0011101101000000" => data <= "100110";
				when "0011101101000001" => data <= "111111";
				when "0011101101000110" => data <= "111111";
				when "0011101101000111" => data <= "111111";
				when "0011101101001000" => data <= "010110";
				when "0011101101001001" => data <= "010110";
				when "0011101101001010" => data <= "100111";
				when "0011101101001011" => data <= "100110";
				when "0011101101001100" => data <= "111111";
				when "0011101101001101" => data <= "111111";
				when "0011101101001110" => data <= "111111";
				when "0011101101010110" => data <= "111111";
				when "0011101101010111" => data <= "100111";
				when "0011101101011000" => data <= "100111";
				when "0011101101011001" => data <= "100111";
				when "0011101101011010" => data <= "100110";
				when "0011101101011011" => data <= "111111";
				when "0011101101101001" => data <= "111111";
				when "0011101101101010" => data <= "100110";
				when "0011101101101011" => data <= "100111";
				when "0011101101101100" => data <= "100111";
				when "0011101101101101" => data <= "100111";
				when "0011101101101110" => data <= "111111";
				when "0011101101110010" => data <= "111111";
				when "0011101101110011" => data <= "100110";
				when "0011101101110100" => data <= "100110";
				when "0011101101110101" => data <= "111111";
				when "0011101101110110" => data <= "111111";
				when "0011110000100111" => data <= "111111";
				when "0011110000101000" => data <= "010010";
				when "0011110000101001" => data <= "010010";
				when "0011110000101010" => data <= "111111";
				when "0011110000101011" => data <= "111111";
				when "0011110000110001" => data <= "111111";
				when "0011110000110010" => data <= "010010";
				when "0011110000110011" => data <= "010010";
				when "0011110000110100" => data <= "111111";
				when "0011110000110101" => data <= "111111";
				when "0011110000111100" => data <= "111111";
				when "0011110000111101" => data <= "111111";
				when "0011110000111110" => data <= "010010";
				when "0011110000111111" => data <= "010010";
				when "0011110001000000" => data <= "010010";
				when "0011110001000001" => data <= "010010";
				when "0011110001000010" => data <= "111111";
				when "0011110001000110" => data <= "111111";
				when "0011110001000111" => data <= "010010";
				when "0011110001001000" => data <= "010010";
				when "0011110001001001" => data <= "010010";
				when "0011110001001010" => data <= "010010";
				when "0011110001001011" => data <= "010110";
				when "0011110001001100" => data <= "111111";
				when "0011110001010110" => data <= "111111";
				when "0011110001010111" => data <= "010111";
				when "0011110001011000" => data <= "010111";
				when "0011110001011001" => data <= "100111";
				when "0011110001011010" => data <= "100111";
				when "0011110001011011" => data <= "111111";
				when "0011110001011100" => data <= "111111";
				when "0011110001011101" => data <= "111111";
				when "0011110001011110" => data <= "111111";
				when "0011110001011111" => data <= "111111";
				when "0011110001100000" => data <= "111111";
				when "0011110001100001" => data <= "111111";
				when "0011110001100010" => data <= "111111";
				when "0011110001101001" => data <= "111111";
				when "0011110001101010" => data <= "010010";
				when "0011110001101011" => data <= "010011";
				when "0011110001101100" => data <= "010011";
				when "0011110001101101" => data <= "010010";
				when "0011110001101110" => data <= "111111";
				when "0011110001101111" => data <= "111111";
				when "0011110001110000" => data <= "111111";
				when "0011110001110001" => data <= "111111";
				when "0011110001110010" => data <= "111111";
				when "0011110001110011" => data <= "010010";
				when "0011110001110100" => data <= "010010";
				when "0011110001110101" => data <= "111111";
				when "0011110001110110" => data <= "111111";
				when "0011110100100111" => data <= "111111";
				when "0011110100101000" => data <= "010010";
				when "0011110100101001" => data <= "010010";
				when "0011110100101010" => data <= "111111";
				when "0011110100101011" => data <= "111111";
				when "0011110100110001" => data <= "111111";
				when "0011110100110010" => data <= "010010";
				when "0011110100110011" => data <= "010010";
				when "0011110100110100" => data <= "111111";
				when "0011110100110101" => data <= "111111";
				when "0011110100111101" => data <= "111111";
				when "0011110100111110" => data <= "111111";
				when "0011110100111111" => data <= "111111";
				when "0011110101000000" => data <= "010010";
				when "0011110101000001" => data <= "010010";
				when "0011110101000010" => data <= "010010";
				when "0011110101000011" => data <= "111111";
				when "0011110101000100" => data <= "111111";
				when "0011110101000101" => data <= "111111";
				when "0011110101000110" => data <= "111111";
				when "0011110101000111" => data <= "010010";
				when "0011110101001000" => data <= "010010";
				when "0011110101001001" => data <= "010010";
				when "0011110101001010" => data <= "010010";
				when "0011110101001011" => data <= "111111";
				when "0011110101010110" => data <= "111111";
				when "0011110101010111" => data <= "010010";
				when "0011110101011000" => data <= "010010";
				when "0011110101011001" => data <= "010011";
				when "0011110101011010" => data <= "010010";
				when "0011110101011011" => data <= "010010";
				when "0011110101011100" => data <= "010010";
				when "0011110101011101" => data <= "010010";
				when "0011110101011110" => data <= "010110";
				when "0011110101011111" => data <= "010110";
				when "0011110101100000" => data <= "010110";
				when "0011110101100001" => data <= "010101";
				when "0011110101100010" => data <= "010101";
				when "0011110101100011" => data <= "111111";
				when "0011110101101001" => data <= "111111";
				when "0011110101101010" => data <= "010010";
				when "0011110101101011" => data <= "010010";
				when "0011110101101100" => data <= "010010";
				when "0011110101101101" => data <= "010011";
				when "0011110101101110" => data <= "010010";
				when "0011110101101111" => data <= "010010";
				when "0011110101110000" => data <= "010110";
				when "0011110101110001" => data <= "010110";
				when "0011110101110010" => data <= "010110";
				when "0011110101110011" => data <= "010010";
				when "0011110101110100" => data <= "111111";
				when "0011111000100111" => data <= "111111";
				when "0011111000101000" => data <= "010010";
				when "0011111000101001" => data <= "010010";
				when "0011111000101010" => data <= "111111";
				when "0011111000101011" => data <= "111111";
				when "0011111000110001" => data <= "111111";
				when "0011111000110010" => data <= "010010";
				when "0011111000110011" => data <= "010010";
				when "0011111000110100" => data <= "111111";
				when "0011111000110101" => data <= "111111";
				when "0011111000111110" => data <= "111111";
				when "0011111000111111" => data <= "111111";
				when "0011111001000000" => data <= "010110";
				when "0011111001000001" => data <= "010010";
				when "0011111001000010" => data <= "010011";
				when "0011111001000011" => data <= "010010";
				when "0011111001000100" => data <= "010010";
				when "0011111001000101" => data <= "111111";
				when "0011111001000110" => data <= "010010";
				when "0011111001000111" => data <= "010011";
				when "0011111001001000" => data <= "010010";
				when "0011111001001001" => data <= "010010";
				when "0011111001001010" => data <= "010010";
				when "0011111001001011" => data <= "111111";
				when "0011111001010110" => data <= "111111";
				when "0011111001010111" => data <= "010010";
				when "0011111001011000" => data <= "010010";
				when "0011111001011001" => data <= "010011";
				when "0011111001011010" => data <= "010010";
				when "0011111001011011" => data <= "010010";
				when "0011111001011100" => data <= "010010";
				when "0011111001011101" => data <= "010010";
				when "0011111001011110" => data <= "010110";
				when "0011111001011111" => data <= "010110";
				when "0011111001100000" => data <= "010110";
				when "0011111001100001" => data <= "010110";
				when "0011111001100010" => data <= "010110";
				when "0011111001100011" => data <= "111111";
				when "0011111001101001" => data <= "111111";
				when "0011111001101010" => data <= "010010";
				when "0011111001101011" => data <= "010010";
				when "0011111001101100" => data <= "010010";
				when "0011111001101101" => data <= "010010";
				when "0011111001101110" => data <= "010010";
				when "0011111001101111" => data <= "010110";
				when "0011111001110000" => data <= "010110";
				when "0011111001110001" => data <= "010110";
				when "0011111001110010" => data <= "010010";
				when "0011111001110011" => data <= "010011";
				when "0011111001110100" => data <= "010010";
				when "0011111001110101" => data <= "111111";
				when "0011111001110110" => data <= "111111";
				when "0011111100100111" => data <= "111111";
				when "0011111100101000" => data <= "010010";
				when "0011111100101001" => data <= "010010";
				when "0011111100101010" => data <= "111111";
				when "0011111100101011" => data <= "111111";
				when "0011111100110001" => data <= "111111";
				when "0011111100110010" => data <= "010010";
				when "0011111100110011" => data <= "010010";
				when "0011111100110100" => data <= "111111";
				when "0011111100110101" => data <= "111111";
				when "0011111100111110" => data <= "111111";
				when "0011111100111111" => data <= "111111";
				when "0011111101000000" => data <= "010110";
				when "0011111101000001" => data <= "010010";
				when "0011111101000010" => data <= "010011";
				when "0011111101000011" => data <= "010010";
				when "0011111101000100" => data <= "010010";
				when "0011111101000101" => data <= "111111";
				when "0011111101000110" => data <= "010010";
				when "0011111101000111" => data <= "010011";
				when "0011111101001000" => data <= "010010";
				when "0011111101001001" => data <= "010010";
				when "0011111101001010" => data <= "010010";
				when "0011111101001011" => data <= "111111";
				when "0011111101010110" => data <= "111111";
				when "0011111101010111" => data <= "010010";
				when "0011111101011000" => data <= "010010";
				when "0011111101011001" => data <= "010011";
				when "0011111101011010" => data <= "010010";
				when "0011111101011011" => data <= "010010";
				when "0011111101011100" => data <= "010010";
				when "0011111101011101" => data <= "010010";
				when "0011111101011110" => data <= "010110";
				when "0011111101011111" => data <= "010110";
				when "0011111101100000" => data <= "010110";
				when "0011111101100001" => data <= "010110";
				when "0011111101100010" => data <= "010110";
				when "0011111101100011" => data <= "111111";
				when "0011111101101001" => data <= "111111";
				when "0011111101101010" => data <= "010010";
				when "0011111101101011" => data <= "010010";
				when "0011111101101100" => data <= "010010";
				when "0011111101101101" => data <= "010010";
				when "0011111101101110" => data <= "010010";
				when "0011111101101111" => data <= "010110";
				when "0011111101110000" => data <= "010110";
				when "0011111101110001" => data <= "010110";
				when "0011111101110010" => data <= "010010";
				when "0011111101110011" => data <= "010011";
				when "0011111101110100" => data <= "010010";
				when "0011111101110101" => data <= "111111";
				when "0011111101110110" => data <= "111111";
				when "0100000000100111" => data <= "111111";
				when "0100000000101000" => data <= "010010";
				when "0100000000101001" => data <= "010010";
				when "0100000000101010" => data <= "111111";
				when "0100000000101011" => data <= "111111";
				when "0100000000110001" => data <= "111111";
				when "0100000000110010" => data <= "010010";
				when "0100000000110011" => data <= "010010";
				when "0100000000110100" => data <= "111111";
				when "0100000000110101" => data <= "111111";
				when "0100000001000000" => data <= "111111";
				when "0100000001000001" => data <= "010010";
				when "0100000001000010" => data <= "010011";
				when "0100000001000011" => data <= "010010";
				when "0100000001000100" => data <= "010010";
				when "0100000001000101" => data <= "010010";
				when "0100000001000110" => data <= "010011";
				when "0100000001000111" => data <= "010011";
				when "0100000001001000" => data <= "010010";
				when "0100000001001001" => data <= "010010";
				when "0100000001001010" => data <= "111111";
				when "0100000001010110" => data <= "111111";
				when "0100000001010111" => data <= "010010";
				when "0100000001011000" => data <= "010010";
				when "0100000001011001" => data <= "010011";
				when "0100000001011010" => data <= "010010";
				when "0100000001011011" => data <= "111111";
				when "0100000001011100" => data <= "111111";
				when "0100000001011101" => data <= "111111";
				when "0100000001011110" => data <= "111111";
				when "0100000001011111" => data <= "111111";
				when "0100000001100000" => data <= "111111";
				when "0100000001100001" => data <= "111111";
				when "0100000001100010" => data <= "111111";
				when "0100000001101001" => data <= "111111";
				when "0100000001101010" => data <= "010010";
				when "0100000001101011" => data <= "010010";
				when "0100000001101100" => data <= "010010";
				when "0100000001101101" => data <= "111111";
				when "0100000001101110" => data <= "111111";
				when "0100000001101111" => data <= "111111";
				when "0100000001110000" => data <= "111111";
				when "0100000001110001" => data <= "111111";
				when "0100000001110010" => data <= "111111";
				when "0100000001110011" => data <= "010011";
				when "0100000001110100" => data <= "010010";
				when "0100000001110101" => data <= "111111";
				when "0100000001110110" => data <= "111111";
				when "0100000100100111" => data <= "111111";
				when "0100000100101000" => data <= "010010";
				when "0100000100101001" => data <= "010010";
				when "0100000100101010" => data <= "111111";
				when "0100000100101011" => data <= "111111";
				when "0100000100110001" => data <= "111111";
				when "0100000100110010" => data <= "010010";
				when "0100000100110011" => data <= "010010";
				when "0100000100110100" => data <= "111111";
				when "0100000100110101" => data <= "111111";
				when "0100000101000000" => data <= "111111";
				when "0100000101000001" => data <= "111111";
				when "0100000101000010" => data <= "010010";
				when "0100000101000011" => data <= "010010";
				when "0100000101000100" => data <= "010010";
				when "0100000101000101" => data <= "010010";
				when "0100000101000110" => data <= "010010";
				when "0100000101000111" => data <= "010010";
				when "0100000101001000" => data <= "111111";
				when "0100000101001001" => data <= "111111";
				when "0100000101001010" => data <= "111111";
				when "0100000101010110" => data <= "111111";
				when "0100000101010111" => data <= "010010";
				when "0100000101011000" => data <= "010010";
				when "0100000101011001" => data <= "010011";
				when "0100000101011010" => data <= "010010";
				when "0100000101011011" => data <= "111111";
				when "0100000101101001" => data <= "111111";
				when "0100000101101010" => data <= "010001";
				when "0100000101101011" => data <= "010001";
				when "0100000101101100" => data <= "010001";
				when "0100000101101101" => data <= "111111";
				when "0100000101110010" => data <= "111111";
				when "0100000101110011" => data <= "010010";
				when "0100000101110100" => data <= "010010";
				when "0100000101110101" => data <= "111111";
				when "0100000101110110" => data <= "111111";
				when "0100001000100111" => data <= "111111";
				when "0100001000101000" => data <= "010010";
				when "0100001000101001" => data <= "010010";
				when "0100001000101010" => data <= "111111";
				when "0100001000101011" => data <= "111111";
				when "0100001000110001" => data <= "111111";
				when "0100001000110010" => data <= "010010";
				when "0100001000110011" => data <= "010010";
				when "0100001000110100" => data <= "111111";
				when "0100001000110101" => data <= "111111";
				when "0100001001000001" => data <= "111111";
				when "0100001001000010" => data <= "010001";
				when "0100001001000011" => data <= "010010";
				when "0100001001000100" => data <= "010010";
				when "0100001001000101" => data <= "010010";
				when "0100001001000110" => data <= "010010";
				when "0100001001000111" => data <= "010010";
				when "0100001001001000" => data <= "111111";
				when "0100001001001001" => data <= "111111";
				when "0100001001010110" => data <= "111111";
				when "0100001001010111" => data <= "010010";
				when "0100001001011000" => data <= "010010";
				when "0100001001011001" => data <= "010010";
				when "0100001001011010" => data <= "010010";
				when "0100001001011011" => data <= "111111";
				when "0100001001101001" => data <= "111111";
				when "0100001001101010" => data <= "010001";
				when "0100001001101011" => data <= "010001";
				when "0100001001101100" => data <= "010001";
				when "0100001001101101" => data <= "111111";
				when "0100001001110010" => data <= "111111";
				when "0100001001110011" => data <= "010010";
				when "0100001001110100" => data <= "010010";
				when "0100001001110101" => data <= "111111";
				when "0100001001110110" => data <= "111111";
				when "0100001100100111" => data <= "111111";
				when "0100001100101000" => data <= "010010";
				when "0100001100101001" => data <= "010010";
				when "0100001100101010" => data <= "111111";
				when "0100001100101011" => data <= "111111";
				when "0100001100101100" => data <= "111111";
				when "0100001100101101" => data <= "111111";
				when "0100001100101110" => data <= "111111";
				when "0100001100101111" => data <= "111111";
				when "0100001100110000" => data <= "111111";
				when "0100001100110001" => data <= "111111";
				when "0100001100110010" => data <= "010010";
				when "0100001100110011" => data <= "010010";
				when "0100001100110100" => data <= "111111";
				when "0100001100110101" => data <= "111111";
				when "0100001101000010" => data <= "111111";
				when "0100001101000011" => data <= "010010";
				when "0100001101000100" => data <= "010010";
				when "0100001101000101" => data <= "010010";
				when "0100001101000110" => data <= "010010";
				when "0100001101000111" => data <= "111111";
				when "0100001101010110" => data <= "111111";
				when "0100001101010111" => data <= "010010";
				when "0100001101011000" => data <= "010010";
				when "0100001101011001" => data <= "010010";
				when "0100001101011010" => data <= "010010";
				when "0100001101011011" => data <= "111111";
				when "0100001101101001" => data <= "111111";
				when "0100001101101010" => data <= "000001";
				when "0100001101101011" => data <= "010001";
				when "0100001101101100" => data <= "010001";
				when "0100001101101101" => data <= "111111";
				when "0100001101110010" => data <= "111111";
				when "0100001101110011" => data <= "010010";
				when "0100001101110100" => data <= "010010";
				when "0100001101110101" => data <= "111111";
				when "0100001101110110" => data <= "111111";
				when "0100010000100111" => data <= "111111";
				when "0100010000101000" => data <= "010010";
				when "0100010000101001" => data <= "010010";
				when "0100010000101010" => data <= "111111";
				when "0100010000101011" => data <= "111111";
				when "0100010000101100" => data <= "111111";
				when "0100010000101101" => data <= "111111";
				when "0100010000101110" => data <= "111111";
				when "0100010000101111" => data <= "111111";
				when "0100010000110000" => data <= "111111";
				when "0100010000110001" => data <= "111111";
				when "0100010000110010" => data <= "010010";
				when "0100010000110011" => data <= "010010";
				when "0100010000110100" => data <= "111111";
				when "0100010000110101" => data <= "111111";
				when "0100010001000010" => data <= "111111";
				when "0100010001000011" => data <= "010010";
				when "0100010001000100" => data <= "010010";
				when "0100010001000101" => data <= "010010";
				when "0100010001000110" => data <= "010010";
				when "0100010001000111" => data <= "111111";
				when "0100010001010110" => data <= "111111";
				when "0100010001010111" => data <= "010010";
				when "0100010001011000" => data <= "010010";
				when "0100010001011001" => data <= "010010";
				when "0100010001011010" => data <= "010010";
				when "0100010001011011" => data <= "111111";
				when "0100010001101001" => data <= "111111";
				when "0100010001101010" => data <= "000001";
				when "0100010001101011" => data <= "010001";
				when "0100010001101100" => data <= "010001";
				when "0100010001101101" => data <= "111111";
				when "0100010001110010" => data <= "111111";
				when "0100010001110011" => data <= "010010";
				when "0100010001110100" => data <= "010010";
				when "0100010001110101" => data <= "111111";
				when "0100010001110110" => data <= "111111";
				when "0100010100100111" => data <= "111111";
				when "0100010100101000" => data <= "010010";
				when "0100010100101001" => data <= "010010";
				when "0100010100101010" => data <= "010001";
				when "0100010100101011" => data <= "010001";
				when "0100010100101100" => data <= "000001";
				when "0100010100101101" => data <= "000001";
				when "0100010100101110" => data <= "010001";
				when "0100010100101111" => data <= "000001";
				when "0100010100110000" => data <= "000001";
				when "0100010100110001" => data <= "010001";
				when "0100010100110010" => data <= "010010";
				when "0100010100110011" => data <= "010010";
				when "0100010100110100" => data <= "111111";
				when "0100010100110101" => data <= "111111";
				when "0100010101000010" => data <= "111111";
				when "0100010101000011" => data <= "000001";
				when "0100010101000100" => data <= "000001";
				when "0100010101000101" => data <= "010010";
				when "0100010101000110" => data <= "010001";
				when "0100010101000111" => data <= "111111";
				when "0100010101010110" => data <= "111111";
				when "0100010101010111" => data <= "010010";
				when "0100010101011000" => data <= "010010";
				when "0100010101011001" => data <= "010010";
				when "0100010101011010" => data <= "010010";
				when "0100010101011011" => data <= "111111";
				when "0100010101011100" => data <= "111111";
				when "0100010101011101" => data <= "111111";
				when "0100010101011110" => data <= "111111";
				when "0100010101011111" => data <= "111111";
				when "0100010101100000" => data <= "111111";
				when "0100010101100001" => data <= "111111";
				when "0100010101100010" => data <= "111111";
				when "0100010101101001" => data <= "111111";
				when "0100010101101010" => data <= "000001";
				when "0100010101101011" => data <= "010001";
				when "0100010101101100" => data <= "010001";
				when "0100010101101101" => data <= "111111";
				when "0100010101110010" => data <= "111111";
				when "0100010101110011" => data <= "010010";
				when "0100010101110100" => data <= "010010";
				when "0100010101110101" => data <= "111111";
				when "0100010101110110" => data <= "111111";
				when "0100011000100111" => data <= "111111";
				when "0100011000101000" => data <= "010001";
				when "0100011000101001" => data <= "010010";
				when "0100011000101010" => data <= "010001";
				when "0100011000101011" => data <= "010001";
				when "0100011000101100" => data <= "000001";
				when "0100011000101101" => data <= "000001";
				when "0100011000101110" => data <= "000001";
				when "0100011000101111" => data <= "000001";
				when "0100011000110000" => data <= "000001";
				when "0100011000110001" => data <= "010001";
				when "0100011000110010" => data <= "010001";
				when "0100011000110011" => data <= "010001";
				when "0100011000110100" => data <= "111111";
				when "0100011000110101" => data <= "111111";
				when "0100011001000011" => data <= "111111";
				when "0100011001000100" => data <= "111111";
				when "0100011001000101" => data <= "010001";
				when "0100011001000110" => data <= "111111";
				when "0100011001010110" => data <= "111111";
				when "0100011001010111" => data <= "000010";
				when "0100011001011000" => data <= "000010";
				when "0100011001011001" => data <= "010010";
				when "0100011001011010" => data <= "010010";
				when "0100011001011011" => data <= "010010";
				when "0100011001011100" => data <= "000010";
				when "0100011001011101" => data <= "000010";
				when "0100011001011110" => data <= "000010";
				when "0100011001011111" => data <= "000010";
				when "0100011001100000" => data <= "010010";
				when "0100011001100001" => data <= "000001";
				when "0100011001100010" => data <= "000001";
				when "0100011001100011" => data <= "111111";
				when "0100011001101001" => data <= "111111";
				when "0100011001101010" => data <= "010001";
				when "0100011001101011" => data <= "010001";
				when "0100011001101100" => data <= "010001";
				when "0100011001101101" => data <= "111111";
				when "0100011001110010" => data <= "111111";
				when "0100011001110011" => data <= "010010";
				when "0100011001110100" => data <= "010010";
				when "0100011001110101" => data <= "111111";
				when "0100011001110110" => data <= "111111";
				when "0100011100101000" => data <= "111111";
				when "0100011100101001" => data <= "111111";
				when "0100011100101010" => data <= "111111";
				when "0100011100101011" => data <= "111111";
				when "0100011100101100" => data <= "111111";
				when "0100011100101101" => data <= "111111";
				when "0100011100101110" => data <= "111111";
				when "0100011100101111" => data <= "111111";
				when "0100011100110000" => data <= "111111";
				when "0100011100110001" => data <= "111111";
				when "0100011100110010" => data <= "111111";
				when "0100011100110011" => data <= "111111";
				when "0100011101000011" => data <= "111111";
				when "0100011101000100" => data <= "111111";
				when "0100011101000101" => data <= "111111";
				when "0100011101000110" => data <= "111111";
				when "0100011101010110" => data <= "111111";
				when "0100011101010111" => data <= "010001";
				when "0100011101011000" => data <= "010001";
				when "0100011101011001" => data <= "000010";
				when "0100011101011010" => data <= "010010";
				when "0100011101011011" => data <= "000010";
				when "0100011101011100" => data <= "010010";
				when "0100011101011101" => data <= "010010";
				when "0100011101011110" => data <= "000010";
				when "0100011101011111" => data <= "000010";
				when "0100011101100000" => data <= "010010";
				when "0100011101100001" => data <= "010001";
				when "0100011101100010" => data <= "010001";
				when "0100011101100011" => data <= "111111";
				when "0100011101101001" => data <= "111111";
				when "0100011101101010" => data <= "010001";
				when "0100011101101011" => data <= "000001";
				when "0100011101101100" => data <= "000001";
				when "0100011101101101" => data <= "111111";
				when "0100011101110010" => data <= "111111";
				when "0100011101110011" => data <= "000001";
				when "0100011101110100" => data <= "000001";
				when "0100011101110101" => data <= "111111";
				when "0100011101110110" => data <= "111111";
				when "0100100001010111" => data <= "111111";
				when "0100100001011000" => data <= "111111";
				when "0100100001011001" => data <= "111111";
				when "0100100001011010" => data <= "111111";
				when "0100100001011011" => data <= "111111";
				when "0100100001011100" => data <= "111111";
				when "0100100001011101" => data <= "111111";
				when "0100100001011110" => data <= "111111";
				when "0100100001011111" => data <= "111111";
				when "0100100001100000" => data <= "111111";
				when "0100100001100001" => data <= "111111";
				when "0100100001100010" => data <= "111111";
				when "0100100001101010" => data <= "111111";
				when "0100100001101011" => data <= "111111";
				when "0100100001101100" => data <= "111111";
				when "0100100001101101" => data <= "111111";
				when "0100100001110011" => data <= "111111";
				when "0100100001110100" => data <= "111111";
				when "0100100101010111" => data <= "111111";
				when "0100100101011000" => data <= "111111";
				when "0100100101011001" => data <= "111111";
				when "0100100101011010" => data <= "111111";
				when "0100100101011011" => data <= "111111";
				when "0100100101011100" => data <= "111111";
				when "0100100101011101" => data <= "111111";
				when "0100100101011110" => data <= "111111";
				when "0100100101011111" => data <= "111111";
				when "0100100101100000" => data <= "111111";
				when "0100100101100001" => data <= "111111";
				when "0100100101100010" => data <= "111111";
				when "0100100101101010" => data <= "111111";
				when "0100100101101011" => data <= "111111";
				when "0100100101101100" => data <= "111111";
				when "0100100101101101" => data <= "111111";
				when "0100100101110011" => data <= "111111";
				when "0100100101110100" => data <= "111111";
				when "0101010000001110" => data <= "111111";
				when "0101010000001111" => data <= "111111";
				when "0101010000010000" => data <= "111111";
				when "0101010000010001" => data <= "111111";
				when "0101010000010010" => data <= "111111";
				when "0101010000010011" => data <= "111111";
				when "0101010000010100" => data <= "111111";
				when "0101010000011001" => data <= "111111";
				when "0101010000011010" => data <= "111111";
				when "0101010000011011" => data <= "111111";
				when "0101010000011100" => data <= "111111";
				when "0101010000011101" => data <= "111111";
				when "0101010000011110" => data <= "111111";
				when "0101010000011111" => data <= "111111";
				when "0101010000100000" => data <= "111111";
				when "0101010000100001" => data <= "111111";
				when "0101010000100111" => data <= "111111";
				when "0101010000101000" => data <= "111111";
				when "0101010000101001" => data <= "111111";
				when "0101010000101010" => data <= "111111";
				when "0101010000101011" => data <= "111111";
				when "0101010000101100" => data <= "111111";
				when "0101010000101101" => data <= "111111";
				when "0101010000110100" => data <= "111111";
				when "0101010000110101" => data <= "111111";
				when "0101010000110110" => data <= "111111";
				when "0101010000110111" => data <= "111111";
				when "0101010000111000" => data <= "111111";
				when "0101010000111001" => data <= "111111";
				when "0101010000111010" => data <= "111111";
				when "0101010001000000" => data <= "111111";
				when "0101010001000001" => data <= "111111";
				when "0101010001000010" => data <= "111111";
				when "0101010001000011" => data <= "111111";
				when "0101010001000100" => data <= "111111";
				when "0101010001000101" => data <= "111111";
				when "0101010001001111" => data <= "111111";
				when "0101010001010000" => data <= "111111";
				when "0101010001010001" => data <= "111111";
				when "0101010001010010" => data <= "111111";
				when "0101010001010011" => data <= "111111";
				when "0101010001010100" => data <= "111111";
				when "0101010001011010" => data <= "111111";
				when "0101010001011011" => data <= "111111";
				when "0101010001011100" => data <= "111111";
				when "0101010001011101" => data <= "111111";
				when "0101010001011110" => data <= "111111";
				when "0101010001011111" => data <= "111111";
				when "0101010001100000" => data <= "111111";
				when "0101010001100110" => data <= "111111";
				when "0101010001100111" => data <= "111111";
				when "0101010001110011" => data <= "111111";
				when "0101010001110100" => data <= "111111";
				when "0101010001110101" => data <= "111111";
				when "0101010001110110" => data <= "111111";
				when "0101010001110111" => data <= "111111";
				when "0101010001111000" => data <= "111111";
				when "0101010001111001" => data <= "111111";
				when "0101010001111111" => data <= "111111";
				when "0101010010000000" => data <= "111111";
				when "0101010010000001" => data <= "111111";
				when "0101010010000010" => data <= "111111";
				when "0101010010000011" => data <= "111111";
				when "0101010010000100" => data <= "111111";
				when "0101010010000101" => data <= "111111";
				when "0101010010001001" => data <= "111111";
				when "0101010010001010" => data <= "111111";
				when "0101010010001011" => data <= "111111";
				when "0101010010001100" => data <= "111111";
				when "0101010010001101" => data <= "111111";
				when "0101010010001110" => data <= "111111";
				when "0101010010001111" => data <= "111111";
				when "0101010010010000" => data <= "111111";
				when "0101010010010001" => data <= "111111";
				when "0101010010010010" => data <= "111111";
				when "0101010100001100" => data <= "111111";
				when "0101010100001101" => data <= "111111";
				when "0101010100001110" => data <= "111111";
				when "0101010100001111" => data <= "111111";
				when "0101010100010000" => data <= "111111";
				when "0101010100010001" => data <= "111111";
				when "0101010100010010" => data <= "111111";
				when "0101010100010011" => data <= "111111";
				when "0101010100010100" => data <= "111111";
				when "0101010100010101" => data <= "111111";
				when "0101010100011001" => data <= "111111";
				when "0101010100011010" => data <= "111111";
				when "0101010100011011" => data <= "111111";
				when "0101010100011100" => data <= "111111";
				when "0101010100011101" => data <= "111111";
				when "0101010100011110" => data <= "111111";
				when "0101010100011111" => data <= "111111";
				when "0101010100100000" => data <= "111111";
				when "0101010100100001" => data <= "111111";
				when "0101010100100010" => data <= "111111";
				when "0101010100100101" => data <= "111111";
				when "0101010100100110" => data <= "111111";
				when "0101010100100111" => data <= "111111";
				when "0101010100101000" => data <= "111111";
				when "0101010100101001" => data <= "111111";
				when "0101010100101010" => data <= "111111";
				when "0101010100101011" => data <= "111111";
				when "0101010100101100" => data <= "111111";
				when "0101010100101101" => data <= "111111";
				when "0101010100101110" => data <= "111111";
				when "0101010100110011" => data <= "111111";
				when "0101010100110100" => data <= "111111";
				when "0101010100110101" => data <= "111111";
				when "0101010100110110" => data <= "111111";
				when "0101010100110111" => data <= "111111";
				when "0101010100111000" => data <= "111111";
				when "0101010100111001" => data <= "111111";
				when "0101010100111010" => data <= "111111";
				when "0101010100111110" => data <= "111111";
				when "0101010100111111" => data <= "111111";
				when "0101010101000000" => data <= "111111";
				when "0101010101000001" => data <= "111111";
				when "0101010101000010" => data <= "111111";
				when "0101010101000011" => data <= "111111";
				when "0101010101000100" => data <= "111111";
				when "0101010101000101" => data <= "111111";
				when "0101010101001101" => data <= "111111";
				when "0101010101001110" => data <= "111111";
				when "0101010101001111" => data <= "111111";
				when "0101010101010000" => data <= "111111";
				when "0101010101010001" => data <= "111111";
				when "0101010101010010" => data <= "111111";
				when "0101010101010011" => data <= "111111";
				when "0101010101010100" => data <= "111111";
				when "0101010101011001" => data <= "111111";
				when "0101010101011010" => data <= "111111";
				when "0101010101011011" => data <= "111111";
				when "0101010101011100" => data <= "111111";
				when "0101010101011101" => data <= "111111";
				when "0101010101011110" => data <= "111111";
				when "0101010101011111" => data <= "111111";
				when "0101010101100000" => data <= "111111";
				when "0101010101100001" => data <= "111111";
				when "0101010101100010" => data <= "111111";
				when "0101010101100110" => data <= "111111";
				when "0101010101100111" => data <= "111111";
				when "0101010101101000" => data <= "111111";
				when "0101010101110010" => data <= "111111";
				when "0101010101110011" => data <= "111111";
				when "0101010101110100" => data <= "111111";
				when "0101010101110101" => data <= "111111";
				when "0101010101110110" => data <= "111111";
				when "0101010101110111" => data <= "111111";
				when "0101010101111000" => data <= "111111";
				when "0101010101111001" => data <= "111111";
				when "0101010101111010" => data <= "111111";
				when "0101010101111011" => data <= "111111";
				when "0101010101111110" => data <= "111111";
				when "0101010101111111" => data <= "111111";
				when "0101010110000000" => data <= "111111";
				when "0101010110000001" => data <= "111111";
				when "0101010110000010" => data <= "111111";
				when "0101010110000011" => data <= "111111";
				when "0101010110000100" => data <= "111111";
				when "0101010110000101" => data <= "111111";
				when "0101010110001000" => data <= "111111";
				when "0101010110001001" => data <= "111111";
				when "0101010110001010" => data <= "111111";
				when "0101010110001011" => data <= "111111";
				when "0101010110001100" => data <= "111111";
				when "0101010110001101" => data <= "111111";
				when "0101010110001110" => data <= "111111";
				when "0101010110001111" => data <= "111111";
				when "0101010110010000" => data <= "111111";
				when "0101010110010001" => data <= "111111";
				when "0101010110010010" => data <= "111111";
				when "0101010110010011" => data <= "111111";
				when "0101010110010100" => data <= "111111";
				when "0101011000001100" => data <= "111111";
				when "0101011000001101" => data <= "111111";
				when "0101011000001110" => data <= "111111";
				when "0101011000010100" => data <= "111111";
				when "0101011000010101" => data <= "111111";
				when "0101011000011001" => data <= "111111";
				when "0101011000011010" => data <= "111111";
				when "0101011000100000" => data <= "111111";
				when "0101011000100001" => data <= "111111";
				when "0101011000100010" => data <= "111111";
				when "0101011000100101" => data <= "111111";
				when "0101011000100110" => data <= "111111";
				when "0101011000100111" => data <= "111111";
				when "0101011000110011" => data <= "111111";
				when "0101011000110100" => data <= "111111";
				when "0101011000110101" => data <= "111111";
				when "0101011000111110" => data <= "111111";
				when "0101011000111111" => data <= "111111";
				when "0101011001000000" => data <= "111111";
				when "0101011001001101" => data <= "111111";
				when "0101011001001110" => data <= "111111";
				when "0101011001001111" => data <= "111111";
				when "0101011001011001" => data <= "111111";
				when "0101011001011010" => data <= "111111";
				when "0101011001100110" => data <= "111111";
				when "0101011001100111" => data <= "111111";
				when "0101011001101000" => data <= "111111";
				when "0101011001110010" => data <= "111111";
				when "0101011001110011" => data <= "111111";
				when "0101011001111110" => data <= "111111";
				when "0101011001111111" => data <= "111111";
				when "0101011010000000" => data <= "111111";
				when "0101011010001101" => data <= "111111";
				when "0101011010001110" => data <= "111111";
				when "0101011010001111" => data <= "111111";
				when "0101011100001100" => data <= "111111";
				when "0101011100001101" => data <= "111111";
				when "0101011100001110" => data <= "111111";
				when "0101011100010100" => data <= "111111";
				when "0101011100010101" => data <= "111111";
				when "0101011100011001" => data <= "111111";
				when "0101011100011010" => data <= "111111";
				when "0101011100100000" => data <= "111111";
				when "0101011100100001" => data <= "111111";
				when "0101011100100010" => data <= "111111";
				when "0101011100100101" => data <= "111111";
				when "0101011100100110" => data <= "111111";
				when "0101011100100111" => data <= "111111";
				when "0101011100110011" => data <= "111111";
				when "0101011100110100" => data <= "111111";
				when "0101011100110101" => data <= "111111";
				when "0101011100111110" => data <= "111111";
				when "0101011100111111" => data <= "111111";
				when "0101011101000000" => data <= "111111";
				when "0101011101001101" => data <= "111111";
				when "0101011101001110" => data <= "111111";
				when "0101011101001111" => data <= "111111";
				when "0101011101011001" => data <= "111111";
				when "0101011101011010" => data <= "111111";
				when "0101011101100110" => data <= "111111";
				when "0101011101100111" => data <= "111111";
				when "0101011101101000" => data <= "111111";
				when "0101011101110010" => data <= "111111";
				when "0101011101110011" => data <= "111111";
				when "0101011101111110" => data <= "111111";
				when "0101011101111111" => data <= "111111";
				when "0101011110000000" => data <= "111111";
				when "0101011110001101" => data <= "111111";
				when "0101011110001110" => data <= "111111";
				when "0101011110001111" => data <= "111111";
				when "0101100000001100" => data <= "111111";
				when "0101100000001101" => data <= "111111";
				when "0101100000001110" => data <= "111111";
				when "0101100000010100" => data <= "111111";
				when "0101100000010101" => data <= "111111";
				when "0101100000011001" => data <= "111111";
				when "0101100000011010" => data <= "111111";
				when "0101100000100000" => data <= "111111";
				when "0101100000100001" => data <= "111111";
				when "0101100000100010" => data <= "111111";
				when "0101100000100101" => data <= "111111";
				when "0101100000100110" => data <= "111111";
				when "0101100000100111" => data <= "111111";
				when "0101100000110011" => data <= "111111";
				when "0101100000110100" => data <= "111111";
				when "0101100000110101" => data <= "111111";
				when "0101100000111110" => data <= "111111";
				when "0101100000111111" => data <= "111111";
				when "0101100001000000" => data <= "111111";
				when "0101100001001101" => data <= "111111";
				when "0101100001001110" => data <= "111111";
				when "0101100001001111" => data <= "111111";
				when "0101100001011001" => data <= "111111";
				when "0101100001011010" => data <= "111111";
				when "0101100001100110" => data <= "111111";
				when "0101100001100111" => data <= "111111";
				when "0101100001101000" => data <= "111111";
				when "0101100001110010" => data <= "111111";
				when "0101100001110011" => data <= "111111";
				when "0101100001111110" => data <= "111111";
				when "0101100001111111" => data <= "111111";
				when "0101100010000000" => data <= "111111";
				when "0101100010001101" => data <= "111111";
				when "0101100010001110" => data <= "111111";
				when "0101100010001111" => data <= "111111";
				when "0101100100001100" => data <= "111111";
				when "0101100100001101" => data <= "111111";
				when "0101100100001110" => data <= "111111";
				when "0101100100010100" => data <= "111111";
				when "0101100100010101" => data <= "111111";
				when "0101100100011001" => data <= "111111";
				when "0101100100011010" => data <= "111111";
				when "0101100100100000" => data <= "111111";
				when "0101100100100001" => data <= "111111";
				when "0101100100100010" => data <= "111111";
				when "0101100100100101" => data <= "111111";
				when "0101100100100110" => data <= "111111";
				when "0101100100100111" => data <= "111111";
				when "0101100100110011" => data <= "111111";
				when "0101100100110100" => data <= "111111";
				when "0101100100110101" => data <= "111111";
				when "0101100100111110" => data <= "111111";
				when "0101100100111111" => data <= "111111";
				when "0101100101000000" => data <= "111111";
				when "0101100101001101" => data <= "111111";
				when "0101100101001110" => data <= "111111";
				when "0101100101001111" => data <= "111111";
				when "0101100101011001" => data <= "111111";
				when "0101100101011010" => data <= "111111";
				when "0101100101100110" => data <= "111111";
				when "0101100101100111" => data <= "111111";
				when "0101100101101000" => data <= "111111";
				when "0101100101110010" => data <= "111111";
				when "0101100101110011" => data <= "111111";
				when "0101100101111110" => data <= "111111";
				when "0101100101111111" => data <= "111111";
				when "0101100110000000" => data <= "111111";
				when "0101100110001101" => data <= "111111";
				when "0101100110001110" => data <= "111111";
				when "0101100110001111" => data <= "111111";
				when "0101101000001100" => data <= "111111";
				when "0101101000001101" => data <= "111111";
				when "0101101000001110" => data <= "111111";
				when "0101101000010100" => data <= "111111";
				when "0101101000010101" => data <= "111111";
				when "0101101000011001" => data <= "111111";
				when "0101101000011010" => data <= "111111";
				when "0101101000100000" => data <= "111111";
				when "0101101000100001" => data <= "111111";
				when "0101101000100010" => data <= "111111";
				when "0101101000100101" => data <= "111111";
				when "0101101000100110" => data <= "111111";
				when "0101101000100111" => data <= "111111";
				when "0101101000110011" => data <= "111111";
				when "0101101000110100" => data <= "111111";
				when "0101101000110101" => data <= "111111";
				when "0101101000111110" => data <= "111111";
				when "0101101000111111" => data <= "111111";
				when "0101101001000000" => data <= "111111";
				when "0101101001001101" => data <= "111111";
				when "0101101001001110" => data <= "111111";
				when "0101101001001111" => data <= "111111";
				when "0101101001011001" => data <= "111111";
				when "0101101001011010" => data <= "111111";
				when "0101101001100110" => data <= "111111";
				when "0101101001100111" => data <= "111111";
				when "0101101001101000" => data <= "111111";
				when "0101101001110010" => data <= "111111";
				when "0101101001110011" => data <= "111111";
				when "0101101001111110" => data <= "111111";
				when "0101101001111111" => data <= "111111";
				when "0101101010000000" => data <= "111111";
				when "0101101010001101" => data <= "111111";
				when "0101101010001110" => data <= "111111";
				when "0101101010001111" => data <= "111111";
				when "0101101100001100" => data <= "111111";
				when "0101101100001101" => data <= "111111";
				when "0101101100001110" => data <= "111111";
				when "0101101100001111" => data <= "111111";
				when "0101101100010000" => data <= "111111";
				when "0101101100010001" => data <= "111111";
				when "0101101100010010" => data <= "111111";
				when "0101101100010011" => data <= "111111";
				when "0101101100010100" => data <= "111111";
				when "0101101100010101" => data <= "111111";
				when "0101101100011001" => data <= "111111";
				when "0101101100011010" => data <= "111111";
				when "0101101100011011" => data <= "111111";
				when "0101101100011100" => data <= "111111";
				when "0101101100011101" => data <= "111111";
				when "0101101100011110" => data <= "111111";
				when "0101101100011111" => data <= "111111";
				when "0101101100100000" => data <= "111111";
				when "0101101100100001" => data <= "111111";
				when "0101101100100010" => data <= "111111";
				when "0101101100100101" => data <= "111111";
				when "0101101100100110" => data <= "111111";
				when "0101101100100111" => data <= "111111";
				when "0101101100101000" => data <= "111111";
				when "0101101100101001" => data <= "111111";
				when "0101101100101010" => data <= "111111";
				when "0101101100101011" => data <= "111111";
				when "0101101100101100" => data <= "111111";
				when "0101101100101101" => data <= "111111";
				when "0101101100101110" => data <= "111111";
				when "0101101100110011" => data <= "111111";
				when "0101101100110100" => data <= "111111";
				when "0101101100110101" => data <= "111111";
				when "0101101100110110" => data <= "111111";
				when "0101101100110111" => data <= "111111";
				when "0101101100111000" => data <= "111111";
				when "0101101100111001" => data <= "111111";
				when "0101101100111010" => data <= "111111";
				when "0101101100111110" => data <= "111111";
				when "0101101100111111" => data <= "111111";
				when "0101101101000000" => data <= "111111";
				when "0101101101000001" => data <= "111111";
				when "0101101101000010" => data <= "111111";
				when "0101101101000011" => data <= "111111";
				when "0101101101000100" => data <= "111111";
				when "0101101101000101" => data <= "111111";
				when "0101101101001101" => data <= "111111";
				when "0101101101001110" => data <= "111111";
				when "0101101101001111" => data <= "111111";
				when "0101101101010000" => data <= "111111";
				when "0101101101010001" => data <= "111111";
				when "0101101101010010" => data <= "111111";
				when "0101101101010011" => data <= "111111";
				when "0101101101010100" => data <= "111111";
				when "0101101101011001" => data <= "111111";
				when "0101101101011010" => data <= "111111";
				when "0101101101011011" => data <= "111111";
				when "0101101101011100" => data <= "111111";
				when "0101101101011101" => data <= "111111";
				when "0101101101011110" => data <= "111111";
				when "0101101101011111" => data <= "111111";
				when "0101101101100000" => data <= "111111";
				when "0101101101100001" => data <= "111111";
				when "0101101101100010" => data <= "111111";
				when "0101101101100110" => data <= "111111";
				when "0101101101100111" => data <= "111111";
				when "0101101101101000" => data <= "111111";
				when "0101101101110010" => data <= "111111";
				when "0101101101110011" => data <= "111111";
				when "0101101101110100" => data <= "111111";
				when "0101101101110101" => data <= "111111";
				when "0101101101110110" => data <= "111111";
				when "0101101101110111" => data <= "111111";
				when "0101101101111000" => data <= "111111";
				when "0101101101111001" => data <= "111111";
				when "0101101101111010" => data <= "111111";
				when "0101101101111011" => data <= "111111";
				when "0101101101111110" => data <= "111111";
				when "0101101101111111" => data <= "111111";
				when "0101101110000000" => data <= "111111";
				when "0101101110001101" => data <= "111111";
				when "0101101110001110" => data <= "111111";
				when "0101101110001111" => data <= "111111";
				when "0101110000001100" => data <= "111111";
				when "0101110000001101" => data <= "111111";
				when "0101110000001110" => data <= "111111";
				when "0101110000001111" => data <= "111111";
				when "0101110000010000" => data <= "111111";
				when "0101110000010001" => data <= "111111";
				when "0101110000010010" => data <= "111111";
				when "0101110000010011" => data <= "111111";
				when "0101110000010100" => data <= "111111";
				when "0101110000011001" => data <= "111111";
				when "0101110000011010" => data <= "111111";
				when "0101110000011011" => data <= "111111";
				when "0101110000011100" => data <= "111111";
				when "0101110000011101" => data <= "111111";
				when "0101110000011110" => data <= "111111";
				when "0101110000011111" => data <= "111111";
				when "0101110000100000" => data <= "111111";
				when "0101110000100001" => data <= "111111";
				when "0101110000100101" => data <= "111111";
				when "0101110000100110" => data <= "111111";
				when "0101110000100111" => data <= "111111";
				when "0101110000101000" => data <= "111111";
				when "0101110000101001" => data <= "111111";
				when "0101110000101010" => data <= "111111";
				when "0101110000101011" => data <= "111111";
				when "0101110000101100" => data <= "111111";
				when "0101110000101101" => data <= "111111";
				when "0101110000101110" => data <= "111111";
				when "0101110000110011" => data <= "111111";
				when "0101110000110100" => data <= "111111";
				when "0101110000110101" => data <= "111111";
				when "0101110000110110" => data <= "111111";
				when "0101110000110111" => data <= "111111";
				when "0101110000111000" => data <= "111111";
				when "0101110000111001" => data <= "111111";
				when "0101110000111010" => data <= "111111";
				when "0101110000111011" => data <= "111111";
				when "0101110001000000" => data <= "111111";
				when "0101110001000001" => data <= "111111";
				when "0101110001000010" => data <= "111111";
				when "0101110001000011" => data <= "111111";
				when "0101110001000100" => data <= "111111";
				when "0101110001000101" => data <= "111111";
				when "0101110001000110" => data <= "111111";
				when "0101110001001111" => data <= "111111";
				when "0101110001010000" => data <= "111111";
				when "0101110001010001" => data <= "111111";
				when "0101110001010010" => data <= "111111";
				when "0101110001010011" => data <= "111111";
				when "0101110001010100" => data <= "111111";
				when "0101110001010101" => data <= "111111";
				when "0101110001011001" => data <= "111111";
				when "0101110001011010" => data <= "111111";
				when "0101110001011011" => data <= "111111";
				when "0101110001011100" => data <= "111111";
				when "0101110001011101" => data <= "111111";
				when "0101110001011110" => data <= "111111";
				when "0101110001011111" => data <= "111111";
				when "0101110001100000" => data <= "111111";
				when "0101110001100001" => data <= "111111";
				when "0101110001100010" => data <= "111111";
				when "0101110001100110" => data <= "111111";
				when "0101110001100111" => data <= "111111";
				when "0101110001101000" => data <= "111111";
				when "0101110001110010" => data <= "111111";
				when "0101110001110011" => data <= "111111";
				when "0101110001110100" => data <= "111111";
				when "0101110001110101" => data <= "111111";
				when "0101110001110110" => data <= "111111";
				when "0101110001110111" => data <= "111111";
				when "0101110001111000" => data <= "111111";
				when "0101110001111001" => data <= "111111";
				when "0101110001111010" => data <= "111111";
				when "0101110001111011" => data <= "111111";
				when "0101110001111110" => data <= "111111";
				when "0101110001111111" => data <= "111111";
				when "0101110010000000" => data <= "111111";
				when "0101110010001101" => data <= "111111";
				when "0101110010001110" => data <= "111111";
				when "0101110010001111" => data <= "111111";
				when "0101110100001100" => data <= "111111";
				when "0101110100001101" => data <= "111111";
				when "0101110100001110" => data <= "111111";
				when "0101110100001111" => data <= "111111";
				when "0101110100010000" => data <= "111111";
				when "0101110100010001" => data <= "111111";
				when "0101110100010010" => data <= "111111";
				when "0101110100010011" => data <= "111111";
				when "0101110100010100" => data <= "111111";
				when "0101110100011001" => data <= "111111";
				when "0101110100011010" => data <= "111111";
				when "0101110100011011" => data <= "111111";
				when "0101110100011100" => data <= "111111";
				when "0101110100011101" => data <= "111111";
				when "0101110100011110" => data <= "111111";
				when "0101110100011111" => data <= "111111";
				when "0101110100100000" => data <= "111111";
				when "0101110100100001" => data <= "111111";
				when "0101110100100101" => data <= "111111";
				when "0101110100100110" => data <= "111111";
				when "0101110100100111" => data <= "111111";
				when "0101110100101000" => data <= "111111";
				when "0101110100101001" => data <= "111111";
				when "0101110100101010" => data <= "111111";
				when "0101110100101011" => data <= "111111";
				when "0101110100101100" => data <= "111111";
				when "0101110100101101" => data <= "111111";
				when "0101110100101110" => data <= "111111";
				when "0101110100110011" => data <= "111111";
				when "0101110100110100" => data <= "111111";
				when "0101110100110101" => data <= "111111";
				when "0101110100110110" => data <= "111111";
				when "0101110100110111" => data <= "111111";
				when "0101110100111000" => data <= "111111";
				when "0101110100111001" => data <= "111111";
				when "0101110100111010" => data <= "111111";
				when "0101110100111011" => data <= "111111";
				when "0101110101000000" => data <= "111111";
				when "0101110101000001" => data <= "111111";
				when "0101110101000010" => data <= "111111";
				when "0101110101000011" => data <= "111111";
				when "0101110101000100" => data <= "111111";
				when "0101110101000101" => data <= "111111";
				when "0101110101000110" => data <= "111111";
				when "0101110101001111" => data <= "111111";
				when "0101110101010000" => data <= "111111";
				when "0101110101010001" => data <= "111111";
				when "0101110101010010" => data <= "111111";
				when "0101110101010011" => data <= "111111";
				when "0101110101010100" => data <= "111111";
				when "0101110101010101" => data <= "111111";
				when "0101110101011001" => data <= "111111";
				when "0101110101011010" => data <= "111111";
				when "0101110101011011" => data <= "111111";
				when "0101110101011100" => data <= "111111";
				when "0101110101011101" => data <= "111111";
				when "0101110101011110" => data <= "111111";
				when "0101110101011111" => data <= "111111";
				when "0101110101100000" => data <= "111111";
				when "0101110101100001" => data <= "111111";
				when "0101110101100010" => data <= "111111";
				when "0101110101100110" => data <= "111111";
				when "0101110101100111" => data <= "111111";
				when "0101110101101000" => data <= "111111";
				when "0101110101110010" => data <= "111111";
				when "0101110101110011" => data <= "111111";
				when "0101110101110100" => data <= "111111";
				when "0101110101110101" => data <= "111111";
				when "0101110101110110" => data <= "111111";
				when "0101110101110111" => data <= "111111";
				when "0101110101111000" => data <= "111111";
				when "0101110101111001" => data <= "111111";
				when "0101110101111010" => data <= "111111";
				when "0101110101111011" => data <= "111111";
				when "0101110101111110" => data <= "111111";
				when "0101110101111111" => data <= "111111";
				when "0101110110000000" => data <= "111111";
				when "0101110110001101" => data <= "111111";
				when "0101110110001110" => data <= "111111";
				when "0101110110001111" => data <= "111111";
				when "0101111000001100" => data <= "111111";
				when "0101111000001101" => data <= "111111";
				when "0101111000001110" => data <= "111111";
				when "0101111000011001" => data <= "111111";
				when "0101111000011010" => data <= "111111";
				when "0101111000100000" => data <= "111111";
				when "0101111000100001" => data <= "111111";
				when "0101111000100010" => data <= "111111";
				when "0101111000100101" => data <= "111111";
				when "0101111000100110" => data <= "111111";
				when "0101111000100111" => data <= "111111";
				when "0101111000111001" => data <= "111111";
				when "0101111000111010" => data <= "111111";
				when "0101111000111011" => data <= "111111";
				when "0101111001000101" => data <= "111111";
				when "0101111001000110" => data <= "111111";
				when "0101111001010100" => data <= "111111";
				when "0101111001010101" => data <= "111111";
				when "0101111001011001" => data <= "111111";
				when "0101111001011010" => data <= "111111";
				when "0101111001100110" => data <= "111111";
				when "0101111001100111" => data <= "111111";
				when "0101111001101000" => data <= "111111";
				when "0101111001110010" => data <= "111111";
				when "0101111001110011" => data <= "111111";
				when "0101111001111110" => data <= "111111";
				when "0101111001111111" => data <= "111111";
				when "0101111010000000" => data <= "111111";
				when "0101111010001101" => data <= "111111";
				when "0101111010001110" => data <= "111111";
				when "0101111010001111" => data <= "111111";
				when "0101111100001100" => data <= "111111";
				when "0101111100001101" => data <= "111111";
				when "0101111100001110" => data <= "111111";
				when "0101111100011001" => data <= "111111";
				when "0101111100011010" => data <= "111111";
				when "0101111100100000" => data <= "111111";
				when "0101111100100001" => data <= "111111";
				when "0101111100100010" => data <= "111111";
				when "0101111100100101" => data <= "111111";
				when "0101111100100110" => data <= "111111";
				when "0101111100100111" => data <= "111111";
				when "0101111100111001" => data <= "111111";
				when "0101111100111010" => data <= "111111";
				when "0101111100111011" => data <= "111111";
				when "0101111101000101" => data <= "111111";
				when "0101111101000110" => data <= "111111";
				when "0101111101010100" => data <= "111111";
				when "0101111101010101" => data <= "111111";
				when "0101111101011001" => data <= "111111";
				when "0101111101011010" => data <= "111111";
				when "0101111101100110" => data <= "111111";
				when "0101111101100111" => data <= "111111";
				when "0101111101101000" => data <= "111111";
				when "0101111101110010" => data <= "111111";
				when "0101111101110011" => data <= "111111";
				when "0101111101111110" => data <= "111111";
				when "0101111101111111" => data <= "111111";
				when "0101111110000000" => data <= "111111";
				when "0101111110001101" => data <= "111111";
				when "0101111110001110" => data <= "111111";
				when "0101111110001111" => data <= "111111";
				when "0110000000001100" => data <= "111111";
				when "0110000000001101" => data <= "111111";
				when "0110000000001110" => data <= "111111";
				when "0110000000011001" => data <= "111111";
				when "0110000000011010" => data <= "111111";
				when "0110000000100000" => data <= "111111";
				when "0110000000100001" => data <= "111111";
				when "0110000000100010" => data <= "111111";
				when "0110000000100101" => data <= "111111";
				when "0110000000100110" => data <= "111111";
				when "0110000000100111" => data <= "111111";
				when "0110000000111001" => data <= "111111";
				when "0110000000111010" => data <= "111111";
				when "0110000000111011" => data <= "111111";
				when "0110000001000101" => data <= "111111";
				when "0110000001000110" => data <= "111111";
				when "0110000001010100" => data <= "111111";
				when "0110000001010101" => data <= "111111";
				when "0110000001011001" => data <= "111111";
				when "0110000001011010" => data <= "111111";
				when "0110000001100110" => data <= "111111";
				when "0110000001100111" => data <= "111111";
				when "0110000001101000" => data <= "111111";
				when "0110000001110010" => data <= "111111";
				when "0110000001110011" => data <= "111111";
				when "0110000001111110" => data <= "111111";
				when "0110000001111111" => data <= "111111";
				when "0110000010000000" => data <= "111111";
				when "0110000010001101" => data <= "111111";
				when "0110000010001110" => data <= "111111";
				when "0110000010001111" => data <= "111111";
				when "0110000100001100" => data <= "111111";
				when "0110000100001101" => data <= "111111";
				when "0110000100001110" => data <= "111111";
				when "0110000100011001" => data <= "111111";
				when "0110000100011010" => data <= "111111";
				when "0110000100100000" => data <= "111111";
				when "0110000100100001" => data <= "111111";
				when "0110000100100010" => data <= "111111";
				when "0110000100100101" => data <= "111111";
				when "0110000100100110" => data <= "111111";
				when "0110000100100111" => data <= "111111";
				when "0110000100111001" => data <= "111111";
				when "0110000100111010" => data <= "111111";
				when "0110000100111011" => data <= "111111";
				when "0110000101000101" => data <= "111111";
				when "0110000101000110" => data <= "111111";
				when "0110000101010100" => data <= "111111";
				when "0110000101010101" => data <= "111111";
				when "0110000101011001" => data <= "111111";
				when "0110000101011010" => data <= "111111";
				when "0110000101100110" => data <= "111111";
				when "0110000101100111" => data <= "111111";
				when "0110000101101000" => data <= "111111";
				when "0110000101110010" => data <= "111111";
				when "0110000101110011" => data <= "111111";
				when "0110000101111110" => data <= "111111";
				when "0110000101111111" => data <= "111111";
				when "0110000110000000" => data <= "111111";
				when "0110000110001101" => data <= "111111";
				when "0110000110001110" => data <= "111111";
				when "0110000110001111" => data <= "111111";
				when "0110001000001100" => data <= "111111";
				when "0110001000001101" => data <= "111111";
				when "0110001000001110" => data <= "111111";
				when "0110001000011001" => data <= "111111";
				when "0110001000011010" => data <= "111111";
				when "0110001000100000" => data <= "111111";
				when "0110001000100001" => data <= "111111";
				when "0110001000100010" => data <= "111111";
				when "0110001000100101" => data <= "111111";
				when "0110001000100110" => data <= "111111";
				when "0110001000100111" => data <= "111111";
				when "0110001000111001" => data <= "111111";
				when "0110001000111010" => data <= "111111";
				when "0110001000111011" => data <= "111111";
				when "0110001001000101" => data <= "111111";
				when "0110001001000110" => data <= "111111";
				when "0110001001010100" => data <= "111111";
				when "0110001001010101" => data <= "111111";
				when "0110001001011001" => data <= "111111";
				when "0110001001011010" => data <= "111111";
				when "0110001001100110" => data <= "111111";
				when "0110001001100111" => data <= "111111";
				when "0110001001101000" => data <= "111111";
				when "0110001001110010" => data <= "111111";
				when "0110001001110011" => data <= "111111";
				when "0110001001111110" => data <= "111111";
				when "0110001001111111" => data <= "111111";
				when "0110001010000000" => data <= "111111";
				when "0110001010001101" => data <= "111111";
				when "0110001010001110" => data <= "111111";
				when "0110001010001111" => data <= "111111";
				when "0110001100001100" => data <= "111111";
				when "0110001100001101" => data <= "111111";
				when "0110001100001110" => data <= "111111";
				when "0110001100011001" => data <= "111111";
				when "0110001100011010" => data <= "111111";
				when "0110001100100000" => data <= "111111";
				when "0110001100100001" => data <= "111111";
				when "0110001100100010" => data <= "111111";
				when "0110001100100101" => data <= "111111";
				when "0110001100100110" => data <= "111111";
				when "0110001100100111" => data <= "111111";
				when "0110001100111001" => data <= "111111";
				when "0110001100111010" => data <= "111111";
				when "0110001100111011" => data <= "111111";
				when "0110001101000101" => data <= "111111";
				when "0110001101000110" => data <= "111111";
				when "0110001101010100" => data <= "111111";
				when "0110001101010101" => data <= "111111";
				when "0110001101011001" => data <= "111111";
				when "0110001101011010" => data <= "111111";
				when "0110001101100110" => data <= "111111";
				when "0110001101100111" => data <= "111111";
				when "0110001101101000" => data <= "111111";
				when "0110001101110010" => data <= "111111";
				when "0110001101110011" => data <= "111111";
				when "0110001101111110" => data <= "111111";
				when "0110001101111111" => data <= "111111";
				when "0110001110000000" => data <= "111111";
				when "0110001110001101" => data <= "111111";
				when "0110001110001110" => data <= "111111";
				when "0110001110001111" => data <= "111111";
				when "0110010000001100" => data <= "111111";
				when "0110010000001101" => data <= "111111";
				when "0110010000001110" => data <= "111111";
				when "0110010000011001" => data <= "111111";
				when "0110010000011010" => data <= "111111";
				when "0110010000100000" => data <= "111111";
				when "0110010000100001" => data <= "111111";
				when "0110010000100010" => data <= "111111";
				when "0110010000100101" => data <= "111111";
				when "0110010000100110" => data <= "111111";
				when "0110010000100111" => data <= "111111";
				when "0110010000111001" => data <= "111111";
				when "0110010000111010" => data <= "111111";
				when "0110010000111011" => data <= "111111";
				when "0110010001000101" => data <= "111111";
				when "0110010001000110" => data <= "111111";
				when "0110010001010100" => data <= "111111";
				when "0110010001010101" => data <= "111111";
				when "0110010001011001" => data <= "111111";
				when "0110010001011010" => data <= "111111";
				when "0110010001100110" => data <= "111111";
				when "0110010001100111" => data <= "111111";
				when "0110010001101000" => data <= "111111";
				when "0110010001110010" => data <= "111111";
				when "0110010001110011" => data <= "111111";
				when "0110010001111110" => data <= "111111";
				when "0110010001111111" => data <= "111111";
				when "0110010010000000" => data <= "111111";
				when "0110010010001101" => data <= "111111";
				when "0110010010001110" => data <= "111111";
				when "0110010010001111" => data <= "111111";
				when "0110010100001100" => data <= "111111";
				when "0110010100001101" => data <= "111111";
				when "0110010100001110" => data <= "111111";
				when "0110010100011001" => data <= "111111";
				when "0110010100011010" => data <= "111111";
				when "0110010100100000" => data <= "111111";
				when "0110010100100001" => data <= "111111";
				when "0110010100100010" => data <= "111111";
				when "0110010100100101" => data <= "111111";
				when "0110010100100110" => data <= "111111";
				when "0110010100100111" => data <= "111111";
				when "0110010100101000" => data <= "111111";
				when "0110010100101001" => data <= "111111";
				when "0110010100101010" => data <= "111111";
				when "0110010100101011" => data <= "111111";
				when "0110010100101100" => data <= "111111";
				when "0110010100101101" => data <= "111111";
				when "0110010100101110" => data <= "111111";
				when "0110010100101111" => data <= "111111";
				when "0110010100110000" => data <= "111111";
				when "0110010100110011" => data <= "111111";
				when "0110010100110100" => data <= "111111";
				when "0110010100110101" => data <= "111111";
				when "0110010100110110" => data <= "111111";
				when "0110010100110111" => data <= "111111";
				when "0110010100111000" => data <= "111111";
				when "0110010100111001" => data <= "111111";
				when "0110010100111010" => data <= "111111";
				when "0110010100111011" => data <= "111111";
				when "0110010101000000" => data <= "111111";
				when "0110010101000001" => data <= "111111";
				when "0110010101000010" => data <= "111111";
				when "0110010101000011" => data <= "111111";
				when "0110010101000100" => data <= "111111";
				when "0110010101000101" => data <= "111111";
				when "0110010101000110" => data <= "111111";
				when "0110010101001111" => data <= "111111";
				when "0110010101010000" => data <= "111111";
				when "0110010101010001" => data <= "111111";
				when "0110010101010010" => data <= "111111";
				when "0110010101010011" => data <= "111111";
				when "0110010101010100" => data <= "111111";
				when "0110010101010101" => data <= "111111";
				when "0110010101011001" => data <= "111111";
				when "0110010101011010" => data <= "111111";
				when "0110010101011011" => data <= "111111";
				when "0110010101011100" => data <= "111111";
				when "0110010101011101" => data <= "111111";
				when "0110010101011110" => data <= "111111";
				when "0110010101011111" => data <= "111111";
				when "0110010101100000" => data <= "111111";
				when "0110010101100001" => data <= "111111";
				when "0110010101100010" => data <= "111111";
				when "0110010101100011" => data <= "111111";
				when "0110010101100110" => data <= "111111";
				when "0110010101100111" => data <= "111111";
				when "0110010101101000" => data <= "111111";
				when "0110010101101001" => data <= "111111";
				when "0110010101101010" => data <= "111111";
				when "0110010101101011" => data <= "111111";
				when "0110010101101100" => data <= "111111";
				when "0110010101101101" => data <= "111111";
				when "0110010101110010" => data <= "111111";
				when "0110010101110011" => data <= "111111";
				when "0110010101110100" => data <= "111111";
				when "0110010101110101" => data <= "111111";
				when "0110010101110110" => data <= "111111";
				when "0110010101110111" => data <= "111111";
				when "0110010101111000" => data <= "111111";
				when "0110010101111001" => data <= "111111";
				when "0110010101111010" => data <= "111111";
				when "0110010101111011" => data <= "111111";
				when "0110010101111100" => data <= "111111";
				when "0110010101111110" => data <= "111111";
				when "0110010101111111" => data <= "111111";
				when "0110010110000000" => data <= "111111";
				when "0110010110000001" => data <= "111111";
				when "0110010110000010" => data <= "111111";
				when "0110010110000011" => data <= "111111";
				when "0110010110000100" => data <= "111111";
				when "0110010110000101" => data <= "111111";
				when "0110010110001101" => data <= "111111";
				when "0110010110001110" => data <= "111111";
				when "0110010110001111" => data <= "111111";
				when "0110011000001110" => data <= "111111";
				when "0110011000011010" => data <= "111111";
				when "0110011000100000" => data <= "111111";
				when "0110011000100001" => data <= "111111";
				when "0110011000100111" => data <= "111111";
				when "0110011000101000" => data <= "111111";
				when "0110011000101001" => data <= "111111";
				when "0110011000101010" => data <= "111111";
				when "0110011000101011" => data <= "111111";
				when "0110011000101100" => data <= "111111";
				when "0110011000101101" => data <= "111111";
				when "0110011000101110" => data <= "111111";
				when "0110011000110011" => data <= "111111";
				when "0110011000110100" => data <= "111111";
				when "0110011000110101" => data <= "111111";
				when "0110011000110110" => data <= "111111";
				when "0110011000110111" => data <= "111111";
				when "0110011000111000" => data <= "111111";
				when "0110011000111001" => data <= "111111";
				when "0110011000111010" => data <= "111111";
				when "0110011001000000" => data <= "111111";
				when "0110011001000001" => data <= "111111";
				when "0110011001000010" => data <= "111111";
				when "0110011001000011" => data <= "111111";
				when "0110011001000100" => data <= "111111";
				when "0110011001000101" => data <= "111111";
				when "0110011001001111" => data <= "111111";
				when "0110011001010000" => data <= "111111";
				when "0110011001010001" => data <= "111111";
				when "0110011001010010" => data <= "111111";
				when "0110011001010011" => data <= "111111";
				when "0110011001010100" => data <= "111111";
				when "0110011001011010" => data <= "111111";
				when "0110011001011011" => data <= "111111";
				when "0110011001011100" => data <= "111111";
				when "0110011001011101" => data <= "111111";
				when "0110011001011110" => data <= "111111";
				when "0110011001011111" => data <= "111111";
				when "0110011001100000" => data <= "111111";
				when "0110011001100001" => data <= "111111";
				when "0110011001100010" => data <= "111111";
				when "0110011001101000" => data <= "111111";
				when "0110011001101001" => data <= "111111";
				when "0110011001101010" => data <= "111111";
				when "0110011001101011" => data <= "111111";
				when "0110011001101100" => data <= "111111";
				when "0110011001101101" => data <= "111111";
				when "0110011001101110" => data <= "111111";
				when "0110011001110011" => data <= "111111";
				when "0110011001110100" => data <= "111111";
				when "0110011001110101" => data <= "111111";
				when "0110011001110110" => data <= "111111";
				when "0110011001110111" => data <= "111111";
				when "0110011001111000" => data <= "111111";
				when "0110011001111001" => data <= "111111";
				when "0110011001111010" => data <= "111111";
				when "0110011001111011" => data <= "111111";
				when "0110011001111111" => data <= "111111";
				when "0110011010000000" => data <= "111111";
				when "0110011010000001" => data <= "111111";
				when "0110011010000010" => data <= "111111";
				when "0110011010000011" => data <= "111111";
				when "0110011010000100" => data <= "111111";
				when "0110011010000101" => data <= "111111";
				when "0110011010001101" => data <= "111111";
				when "0110011010001110" => data <= "111111";
				when "0110011010001111" => data <= "111111";
				when "0110011100001110" => data <= "111111";
				when "0110011100011010" => data <= "111111";
				when "0110011100100000" => data <= "111111";
				when "0110011100100001" => data <= "111111";
				when "0110011100100111" => data <= "111111";
				when "0110011100101000" => data <= "111111";
				when "0110011100101001" => data <= "111111";
				when "0110011100101010" => data <= "111111";
				when "0110011100101011" => data <= "111111";
				when "0110011100101100" => data <= "111111";
				when "0110011100101101" => data <= "111111";
				when "0110011100101110" => data <= "111111";
				when "0110011100110011" => data <= "111111";
				when "0110011100110100" => data <= "111111";
				when "0110011100110101" => data <= "111111";
				when "0110011100110110" => data <= "111111";
				when "0110011100110111" => data <= "111111";
				when "0110011100111000" => data <= "111111";
				when "0110011100111001" => data <= "111111";
				when "0110011100111010" => data <= "111111";
				when "0110011101000000" => data <= "111111";
				when "0110011101000001" => data <= "111111";
				when "0110011101000010" => data <= "111111";
				when "0110011101000011" => data <= "111111";
				when "0110011101000100" => data <= "111111";
				when "0110011101000101" => data <= "111111";
				when "0110011101001111" => data <= "111111";
				when "0110011101010000" => data <= "111111";
				when "0110011101010001" => data <= "111111";
				when "0110011101010010" => data <= "111111";
				when "0110011101010011" => data <= "111111";
				when "0110011101010100" => data <= "111111";
				when "0110011101011010" => data <= "111111";
				when "0110011101011011" => data <= "111111";
				when "0110011101011100" => data <= "111111";
				when "0110011101011101" => data <= "111111";
				when "0110011101011110" => data <= "111111";
				when "0110011101011111" => data <= "111111";
				when "0110011101100000" => data <= "111111";
				when "0110011101100001" => data <= "111111";
				when "0110011101100010" => data <= "111111";
				when "0110011101101000" => data <= "111111";
				when "0110011101101001" => data <= "111111";
				when "0110011101101010" => data <= "111111";
				when "0110011101101011" => data <= "111111";
				when "0110011101101100" => data <= "111111";
				when "0110011101101101" => data <= "111111";
				when "0110011101101110" => data <= "111111";
				when "0110011101110011" => data <= "111111";
				when "0110011101110100" => data <= "111111";
				when "0110011101110101" => data <= "111111";
				when "0110011101110110" => data <= "111111";
				when "0110011101110111" => data <= "111111";
				when "0110011101111000" => data <= "111111";
				when "0110011101111001" => data <= "111111";
				when "0110011101111010" => data <= "111111";
				when "0110011101111011" => data <= "111111";
				when "0110011101111111" => data <= "111111";
				when "0110011110000000" => data <= "111111";
				when "0110011110000001" => data <= "111111";
				when "0110011110000010" => data <= "111111";
				when "0110011110000011" => data <= "111111";
				when "0110011110000100" => data <= "111111";
				when "0110011110000101" => data <= "111111";
				when "0110011110001101" => data <= "111111";
				when "0110011110001110" => data <= "111111";
				when "0110011110001111" => data <= "111111";
				when others => data <= "000000";
			end case;
              		end if; 
              	end process; 
              end;